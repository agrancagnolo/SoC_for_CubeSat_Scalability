* NGSPICE file created from Mixer.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_01v8_Y6SADL a_n210_n1149# a_n50_n1063# a_50_n975# a_n108_n975#
X0 a_50_n975# a_n50_n1063# a_n108_n975# a_n210_n1149# sky130_fd_pr__nfet_01v8 ad=2.8275 pd=20.08 as=2.8275 ps=20.08 w=9.75 l=0.5
**devattr s=113100,4016 d=113100,4016
C0 a_50_n975# a_n50_n1063# 0.062988f
C1 a_n108_n975# a_n50_n1063# 0.064897f
C2 a_50_n975# a_n108_n975# 0.336849f
C3 a_50_n975# a_n210_n1149# 0.819905f
C4 a_n108_n975# a_n210_n1149# 0.611795f
C5 a_n50_n1063# a_n210_n1149# 0.48776f
.ends

.subckt sky130_fd_pr__nfet_01v8_Y6FLEL a_n210_n1149# a_n50_n1063# a_50_n975# a_n108_n975#
X0 a_50_n975# a_n50_n1063# a_n108_n975# a_n210_n1149# sky130_fd_pr__nfet_01v8 ad=2.8275 pd=20.08 as=2.8275 ps=20.08 w=9.75 l=0.5
**devattr s=113100,4016 d=113100,4016
C0 a_50_n975# a_n50_n1063# 0.064897f
C1 a_n108_n975# a_n50_n1063# 0.062988f
C2 a_50_n975# a_n108_n975# 0.336849f
C3 a_50_n975# a_n210_n1149# 0.611795f
C4 a_n108_n975# a_n210_n1149# 0.821788f
C5 a_n50_n1063# a_n210_n1149# 0.48776f
.ends

.subckt sky130_fd_pr__nfet_01v8_PZKCVB a_n50_n1038# a_50_n950# a_n108_n950# a_n210_n1124#
X0 a_50_n950# a_n50_n1038# a_n108_n950# a_n210_n1124# sky130_fd_pr__nfet_01v8 ad=2.755 pd=19.58 as=2.755 ps=19.58 w=9.5 l=0.5
**devattr s=110200,3916 d=110200,3916
C0 a_50_n950# a_n50_n1038# 0.063286f
C1 a_n108_n950# a_n50_n1038# 0.109746f
C2 a_50_n950# a_n108_n950# 0.578324f
C3 a_50_n950# a_n210_n1124# 0.783383f
C4 a_n108_n950# a_n210_n1124# 1.06096f
C5 a_n50_n1038# a_n210_n1124# 0.512003f
.ends

.subckt sky130_fd_pr__nfet_01v8_PMG9RB a_n50_n1038# a_50_n950# a_n108_n950# a_n210_n1124#
X0 a_50_n950# a_n50_n1038# a_n108_n950# a_n210_n1124# sky130_fd_pr__nfet_01v8 ad=2.755 pd=19.58 as=2.755 ps=19.58 w=9.5 l=0.5
**devattr s=110200,3916 d=110200,3916
C0 a_50_n950# a_n50_n1038# 0.034295f
C1 a_n108_n950# a_n50_n1038# 0.05164f
C2 a_50_n950# a_n108_n950# 0.418488f
C3 a_50_n950# a_n210_n1124# 0.656996f
C4 a_n108_n950# a_n210_n1124# 0.757556f
C5 a_n50_n1038# a_n210_n1124# 0.518551f
.ends

.subckt sky130_fd_pr__nfet_01v8_8XPPYK a_n123_n1515# a_n65_n1570# a_65_n1515# a_n225_n1689#
X0 a_65_n1515# a_n65_n1570# a_n123_n1515# a_n225_n1689# sky130_fd_pr__nfet_01v8 ad=4.3935 pd=30.88 as=4.3935 ps=30.88 w=15.15 l=0.65
**devattr s=175740,6176 d=175740,6176
C0 a_65_n1515# a_n65_n1570# 0.192222f
C1 a_n123_n1515# a_n65_n1570# 0.192222f
C2 a_65_n1515# a_n123_n1515# 0.909199f
C3 a_65_n1515# a_n225_n1689# 1.32867f
C4 a_n123_n1515# a_n225_n1689# 1.32867f
C5 a_n65_n1570# a_n225_n1689# 0.570216f
.ends

.subckt sky130_fd_pr__nfet_01v8_Z6VF7Q a_n50_n1038# a_50_n950# a_n108_n950# a_n210_n1124#
X0 a_50_n950# a_n50_n1038# a_n108_n950# a_n210_n1124# sky130_fd_pr__nfet_01v8 ad=2.755 pd=19.58 as=2.755 ps=19.58 w=9.5 l=0.5
**devattr s=110200,3916 d=110200,3916
C0 a_50_n950# a_n50_n1038# 0.074932f
C1 a_n108_n950# a_n50_n1038# 0.077286f
C2 a_50_n950# a_n108_n950# 0.576568f
C3 a_50_n950# a_n210_n1124# 0.750751f
C4 a_n108_n950# a_n210_n1124# 0.764718f
C5 a_n50_n1038# a_n210_n1124# 0.48776f
.ends

.subckt sky130_fd_pr__nfet_01v8_Z9V85Y a_n50_n1038# a_50_n950# a_n108_n950# a_n210_n1124#
X0 a_50_n950# a_n50_n1038# a_n108_n950# a_n210_n1124# sky130_fd_pr__nfet_01v8 ad=2.755 pd=19.58 as=2.755 ps=19.58 w=9.5 l=0.5
**devattr s=110200,3916 d=110200,3916
C0 a_50_n950# a_n50_n1038# 0.074932f
C1 a_n108_n950# a_n50_n1038# 0.05164f
C2 a_50_n950# a_n108_n950# 0.420437f
C3 a_50_n950# a_n210_n1124# 0.685981f
C4 a_n108_n950# a_n210_n1124# 0.547951f
C5 a_n50_n1038# a_n210_n1124# 0.48776f
.ends

.subckt sky130_fd_pr__nfet_01v8_VJM6P6 a_n210_n1149# a_n50_n1063# a_50_n975# a_n108_n975#
X0 a_50_n975# a_n50_n1063# a_n108_n975# a_n210_n1149# sky130_fd_pr__nfet_01v8 ad=2.8275 pd=20.08 as=2.8275 ps=20.08 w=9.75 l=0.5
**devattr s=113100,4016 d=113100,4016
C0 a_50_n975# a_n50_n1063# 0.052879f
C1 a_n108_n975# a_n50_n1063# 0.052879f
C2 a_50_n975# a_n108_n975# 0.387039f
C3 a_50_n975# a_n210_n1149# 0.499622f
C4 a_n108_n975# a_n210_n1149# 0.499622f
C5 a_n50_n1063# a_n210_n1149# 0.48776f
.ends

.subckt sky130_fd_pr__nfet_01v8_HQ3Y9H a_n210_n1149# a_n50_n1063# a_50_n975# a_n108_n975#
X0 a_50_n975# a_n50_n1063# a_n108_n975# a_n210_n1149# sky130_fd_pr__nfet_01v8 ad=2.8275 pd=20.08 as=2.8275 ps=20.08 w=9.75 l=0.5
**devattr s=113100,4016 d=113100,4016
C0 a_50_n975# a_n50_n1063# 0.065024f
C1 a_n108_n975# a_n50_n1063# 0.065024f
C2 a_50_n975# a_n108_n975# 0.601683f
C3 a_50_n975# a_n210_n1149# 0.868072f
C4 a_n108_n975# a_n210_n1149# 0.868072f
C5 a_n50_n1063# a_n210_n1149# 0.48776f
.ends

.subckt sky130_fd_pr__pfet_01v8_JCZH34 a_n50_n967# a_n108_n870# w_n246_n1089# a_50_n870#
+ VSUBS
X0 a_50_n870# a_n50_n967# a_n108_n870# w_n246_n1089# sky130_fd_pr__pfet_01v8 ad=2.523 pd=17.98 as=2.523 ps=17.98 w=8.7 l=0.5
**devattr s=100920,3596 d=100920,3596
C0 a_n108_n870# w_n246_n1089# 0.286555f
C1 a_50_n870# w_n246_n1089# 0.286555f
C2 a_n50_n967# w_n246_n1089# 0.315361f
C3 a_50_n870# a_n108_n870# 0.393711f
C4 a_n108_n870# a_n50_n967# 0.05833f
C5 a_50_n870# a_n50_n967# 0.05833f
C6 a_50_n870# VSUBS 0.199473f
C7 a_n108_n870# VSUBS 0.199473f
C8 a_n50_n967# VSUBS 0.187452f
C9 w_n246_n1089# VSUBS 4.63286f
.ends

.subckt sky130_fd_pr__pfet_01v8_9F3ELE a_n50_n297# a_50_n200# a_n108_n200# w_n246_n419#
+ VSUBS
X0 a_50_n200# a_n50_n297# a_n108_n200# w_n246_n419# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
**devattr s=23200,916 d=23200,916
C0 a_n108_n200# w_n246_n419# 0.14569f
C1 a_50_n200# w_n246_n419# 0.147195f
C2 a_n50_n297# w_n246_n419# 0.315117f
C3 a_50_n200# a_n108_n200# 0.094372f
C4 a_n108_n200# a_n50_n297# 0.017016f
C5 a_50_n200# a_n50_n297# 0.017016f
C6 a_50_n200# VSUBS 0.084165f
C7 a_n108_n200# VSUBS 0.0856f
C8 a_n50_n297# VSUBS 0.16872f
C9 w_n246_n419# VSUBS 1.8552f
.ends

.subckt sky130_fd_pr__pfet_01v8_4F365H a_n50_n297# a_50_n200# a_n108_n200# w_n246_n419#
+ VSUBS
X0 a_50_n200# a_n50_n297# a_n108_n200# w_n246_n419# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
**devattr s=23200,916 d=23200,916
C0 a_n108_n200# w_n246_n419# 0.140472f
C1 a_50_n200# w_n246_n419# 0.162983f
C2 a_n50_n297# w_n246_n419# 0.315117f
C3 a_50_n200# a_n108_n200# 0.133283f
C4 a_n108_n200# a_n50_n297# 0.017016f
C5 a_50_n200# a_n50_n297# 0.028662f
C6 a_50_n200# VSUBS 0.11652f
C7 a_n108_n200# VSUBS 0.067516f
C8 a_n50_n297# VSUBS 0.16872f
C9 w_n246_n419# VSUBS 1.85116f
.ends

.subckt sky130_fd_pr__pfet_01v8_53Y4NB a_n50_n967# a_n108_n870# w_n246_n1089# a_50_n870#
+ VSUBS
X0 a_50_n870# a_n50_n967# a_n108_n870# w_n246_n1089# sky130_fd_pr__pfet_01v8 ad=2.523 pd=17.98 as=2.523 ps=17.98 w=8.7 l=0.5
**devattr s=100920,3596 d=100920,3596
C0 a_n108_n870# w_n246_n1089# 0.394773f
C1 a_50_n870# w_n246_n1089# 0.394773f
C2 a_n50_n967# w_n246_n1089# 0.310821f
C3 a_50_n870# a_n108_n870# 0.546531f
C4 a_n108_n870# a_n50_n967# 0.07964f
C5 a_50_n870# a_n50_n967# 0.07964f
C6 a_50_n870# VSUBS 0.277547f
C7 a_n108_n870# VSUBS 0.277547f
C8 a_n50_n967# VSUBS 0.18394f
C9 w_n246_n1089# VSUBS 4.57436f
.ends

.subckt Mixer vdd gnd vlo- out- vlo+ vbias2 vbias3 vrf+ vrf- vtail vbias1 out+
XXM1 gnd vrf+ m1_5180_850# m1_4048_1162# sky130_fd_pr__nfet_01v8_Y6SADL
XXM2 gnd vrf- m1_5180_850# m1_4436_2196# sky130_fd_pr__nfet_01v8_Y6FLEL
XXM3 vlo- m1_962_656# out+ gnd sky130_fd_pr__nfet_01v8_PZKCVB
XXM4 vlo+ m1_962_656# out- gnd sky130_fd_pr__nfet_01v8_PMG9RB
XXMTAIL m1_5180_850# vtail gnd gnd sky130_fd_pr__nfet_01v8_8XPPYK
XXM5 vlo+ m1_2744_894# out+ gnd sky130_fd_pr__nfet_01v8_Z6VF7Q
XXM6 vlo- m1_2744_894# out- gnd sky130_fd_pr__nfet_01v8_Z9V85Y
XXM7 gnd vbias1 m1_4048_1162# m1_962_656# sky130_fd_pr__nfet_01v8_VJM6P6
XXM8 gnd vbias1 m1_4436_2196# m1_2744_894# sky130_fd_pr__nfet_01v8_HQ3Y9H
XXM9 vbias2 out+ vdd vdd gnd sky130_fd_pr__pfet_01v8_JCZH34
XXMci2 vbias3 vdd m1_2744_894# vdd gnd sky130_fd_pr__pfet_01v8_9F3ELE
XXMci1 vbias3 vdd m1_962_656# vdd gnd sky130_fd_pr__pfet_01v8_4F365H
XXM10 vbias2 out- vdd vdd gnd sky130_fd_pr__pfet_01v8_53Y4NB
C0 vbias1 vrf+ 0.04072f
C1 m1_4436_2196# vrf+ 0.090483f
C2 vrf- m1_4436_2196# 0.006232f
C3 m1_4048_1162# m1_2744_894# 0.169109f
C4 m1_4048_1162# m1_5180_850# 0.001308f
C5 vbias1 m1_2744_894# 0.174568f
C6 vdd vbias2 0.653058f
C7 vbias1 m1_5180_850# 0.003178f
C8 m1_2744_894# out- 0.351103f
C9 m1_4436_2196# m1_2744_894# 3.71e-20
C10 vrf- vrf+ 0.092405f
C11 m1_2744_894# vlo+ 0.008106f
C12 m1_4436_2196# m1_5180_850# 0.125253f
C13 out- vdd 0.381582f
C14 m1_4436_2196# vtail 1.8e-19
C15 m1_962_656# m1_4048_1162# 0.02315f
C16 m1_962_656# vbias2 0.006527f
C17 vlo- m1_4048_1162# 1.88e-19
C18 m1_962_656# vbias1 0.041703f
C19 out+ vbias2 0.014007f
C20 vlo- vbias1 0.005311f
C21 m1_962_656# out- 0.764945f
C22 m1_962_656# m1_4436_2196# 0.002144f
C23 m1_962_656# vlo+ 0.251472f
C24 out+ out- 0.47663f
C25 m1_2744_894# vrf+ 6.91e-20
C26 out+ vlo+ 0.36689f
C27 vlo- out- 0.047432f
C28 m1_5180_850# vrf+ 0.002f
C29 vrf- m1_5180_850# 0.12077f
C30 vlo- m1_4436_2196# 7.73e-20
C31 vlo- vlo+ 0.254583f
C32 vtail vrf+ 6.55e-20
C33 vrf- vtail 0.003585f
C34 vbias3 vbias2 2.57e-20
C35 vbias3 out- 0.006336f
C36 m1_962_656# vrf+ 7.65e-19
C37 m1_2744_894# m1_5180_850# 8.59e-19
C38 m1_2744_894# vdd 0.185584f
C39 vtail m1_5180_850# 0.005493f
C40 m1_962_656# m1_2744_894# 0.444609f
C41 m1_962_656# m1_5180_850# 0.011578f
C42 out+ m1_2744_894# 0.001419f
C43 m1_962_656# vdd 0.171392f
C44 vlo- m1_2744_894# 0.057464f
C45 out+ vdd 0.139936f
C46 vbias3 m1_2744_894# 0.109264f
C47 out+ m1_962_656# 0.382396f
C48 vbias3 vdd 0.237773f
C49 vlo- m1_962_656# 0.711116f
C50 vlo- out+ 0.104122f
C51 vbias1 m1_4048_1162# 0.066573f
C52 m1_962_656# vbias3 0.025101f
C53 m1_4048_1162# m1_4436_2196# 0.190177f
C54 out- vbias2 0.08841f
C55 vbias1 out- 1.9e-21
C56 vbias1 vlo+ 6.89e-21
C57 vlo+ out- 0.408377f
C58 m1_4048_1162# vrf+ 0.00113f
C59 vbias3 gnd 0.523372f
C60 vdd gnd 14.571484f
C61 vbias2 gnd 0.365475f
C62 m1_4436_2196# gnd 1.780702f
C63 m1_4048_1162# gnd 1.191069f
C64 vbias1 gnd 1.369267f
C65 m1_2744_894# gnd 3.669666f
C66 vtail gnd 1.028648f
C67 out- gnd 3.201187f
C68 vlo+ gnd 1.790222f
C69 m1_962_656# gnd 4.271135f
C70 out+ gnd 4.04321f
C71 vlo- gnd 2.191175f
C72 vrf- gnd 0.655737f
C73 m1_5180_850# gnd 2.748746f
C74 vrf+ gnd 0.658237f
.ends

