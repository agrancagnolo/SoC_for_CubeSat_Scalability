VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO signal_generator
  CLASS BLOCK ;
  FOREIGN signal_generator ;
  ORIGIN 0.000 0.000 ;
  SIZE 1200.000 BY 1200.000 ;
  PIN io_analog[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 32.680 1200.000 33.280 ;
    END
  END io_analog[0]
  PIN io_analog[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 250.280 1200.000 250.880 ;
    END
  END io_analog[10]
  PIN io_analog[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 54.440 1200.000 55.040 ;
    END
  END io_analog[1]
  PIN io_analog[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 76.200 1200.000 76.800 ;
    END
  END io_analog[2]
  PIN io_analog[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 97.960 1200.000 98.560 ;
    END
  END io_analog[3]
  PIN io_analog[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 119.720 1200.000 120.320 ;
    END
  END io_analog[4]
  PIN io_analog[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 141.480 1200.000 142.080 ;
    END
  END io_analog[5]
  PIN io_analog[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 163.240 1200.000 163.840 ;
    END
  END io_analog[6]
  PIN io_analog[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 185.000 1200.000 185.600 ;
    END
  END io_analog[7]
  PIN io_analog[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1196.000 206.760 1200.000 207.360 ;
    END
  END io_analog[8]
  PIN io_analog[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1196.000 228.520 1200.000 229.120 ;
    END
  END io_analog[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 272.040 1200.000 272.640 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 924.840 1200.000 925.440 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 990.120 1200.000 990.720 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1055.400 1200.000 1056.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1120.680 1200.000 1121.280 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1166.920 4.000 1167.520 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1077.160 4.000 1077.760 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 987.400 4.000 988.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 897.640 4.000 898.240 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 807.880 4.000 808.480 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 718.120 4.000 718.720 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 337.320 1200.000 337.920 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 628.360 4.000 628.960 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 538.600 4.000 539.200 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 448.840 4.000 449.440 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 359.080 4.000 359.680 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 269.320 4.000 269.920 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 179.560 4.000 180.160 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.800 4.000 90.400 ;
    END
  END io_in[26]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 402.600 1200.000 403.200 ;
    END
  END io_in[2]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 467.880 1200.000 468.480 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 533.160 1200.000 533.760 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 598.440 1200.000 599.040 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 663.720 1200.000 664.320 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 729.000 1200.000 729.600 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 794.280 1200.000 794.880 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 859.560 1200.000 860.160 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 315.560 1200.000 316.160 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 968.360 1200.000 968.960 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1033.640 1200.000 1034.240 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1098.920 1200.000 1099.520 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1164.200 1200.000 1164.800 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1107.080 4.000 1107.680 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1017.320 4.000 1017.920 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 927.560 4.000 928.160 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 837.800 4.000 838.400 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 748.040 4.000 748.640 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 658.280 4.000 658.880 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 380.840 1200.000 381.440 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 568.520 4.000 569.120 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 478.760 4.000 479.360 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 389.000 4.000 389.600 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.240 4.000 299.840 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 209.480 4.000 210.080 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.720 4.000 120.320 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.960 4.000 30.560 ;
    END
  END io_oeb[26]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 446.120 1200.000 446.720 ;
    END
  END io_oeb[2]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 511.400 1200.000 512.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 576.680 1200.000 577.280 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 641.960 1200.000 642.560 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 707.240 1200.000 707.840 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 772.520 1200.000 773.120 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 837.800 1200.000 838.400 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 903.080 1200.000 903.680 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 293.800 1200.000 294.400 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 1196.000 946.600 1200.000 947.200 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1011.880 1200.000 1012.480 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1077.160 1200.000 1077.760 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1142.440 1200.000 1143.040 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1137.000 4.000 1137.600 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1047.240 4.000 1047.840 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 957.480 4.000 958.080 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 867.720 4.000 868.320 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 777.960 4.000 778.560 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 688.200 4.000 688.800 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 359.080 1200.000 359.680 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 598.440 4.000 599.040 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 508.680 4.000 509.280 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 418.920 4.000 419.520 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 329.160 4.000 329.760 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 239.400 4.000 240.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.880 4.000 60.480 ;
    END
  END io_out[26]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 424.360 1200.000 424.960 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 489.640 1200.000 490.240 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 554.920 1200.000 555.520 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 620.200 1200.000 620.800 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 685.480 1200.000 686.080 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 1196.000 750.760 1200.000 751.360 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 1196.000 816.040 1200.000 816.640 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 1196.000 881.320 1200.000 881.920 ;
    END
  END io_out[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -4.480 0.880 -1.480 1198.640 ;
    END
    PORT
      LAYER met5 ;
        RECT -4.480 0.880 1204.160 3.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -4.480 1195.640 1204.160 1198.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 1201.160 0.880 1204.160 1198.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 4.520 -3.820 6.520 1203.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 69.520 -3.820 71.520 1203.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 134.520 -3.820 136.520 99.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 134.520 501.440 136.520 549.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 134.520 951.440 136.520 1140.805 ;
    END
    PORT
      LAYER met4 ;
        RECT 134.520 1163.365 136.520 1203.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 199.520 -3.820 201.520 99.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 199.520 501.440 201.520 549.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 199.520 951.440 201.520 1203.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 264.520 -3.820 266.520 99.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 264.520 501.440 266.520 549.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 264.520 951.440 266.520 1203.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 329.520 -3.820 331.520 99.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 329.520 501.440 331.520 549.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 329.520 951.440 331.520 1203.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 394.520 -3.820 396.520 99.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 394.520 501.440 396.520 549.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 394.520 951.440 396.520 1203.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 459.520 -3.820 461.520 99.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 459.520 501.440 461.520 549.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 459.520 951.440 461.520 1136.855 ;
    END
    PORT
      LAYER met4 ;
        RECT 459.520 1159.415 461.520 1203.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 524.520 -3.820 526.520 1203.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 589.520 -3.820 591.520 1203.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 654.520 -3.820 656.520 1203.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 719.520 -3.820 721.520 1203.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 784.520 -3.820 786.520 1203.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 849.520 -3.820 851.520 1203.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 914.520 -3.820 916.520 1203.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 979.520 -3.820 981.520 1203.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1044.520 -3.820 1046.520 1203.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1109.520 -3.820 1111.520 1203.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1174.520 -3.820 1176.520 1203.340 ;
    END
    PORT
      LAYER met5 ;
        RECT -9.180 9.880 1208.860 11.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -9.180 74.880 1208.860 76.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -9.180 139.880 66.420 141.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -9.180 204.880 166.200 206.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -9.180 269.880 166.200 271.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -9.180 334.880 66.420 336.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -9.180 399.880 66.420 401.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -9.180 464.880 66.420 466.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -9.180 529.880 1208.860 531.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -9.180 594.880 66.420 596.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -9.180 659.880 66.420 661.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -9.180 724.880 166.200 726.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -9.180 789.880 166.200 791.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -9.180 854.880 66.420 856.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -9.180 919.880 66.420 921.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -9.180 984.880 1208.860 986.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -9.180 1049.880 1208.860 1051.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -9.180 1114.880 1208.860 1116.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -9.180 1179.880 1208.860 1181.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 353.160 269.880 1208.860 271.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 353.160 724.880 1208.860 726.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 353.160 789.880 1208.860 791.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 396.530 204.880 1208.860 206.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 524.520 139.880 1208.860 141.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 524.520 659.880 1208.860 661.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 524.520 854.880 1208.860 856.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 526.320 334.880 1208.860 336.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 526.320 399.880 1208.860 401.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 526.320 464.880 1208.860 466.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 526.320 594.880 1208.860 596.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 526.320 919.880 1208.860 921.880 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -9.180 -3.820 -6.180 1203.340 ;
    END
    PORT
      LAYER met5 ;
        RECT -9.180 -3.820 1208.860 -0.820 ;
    END
    PORT
      LAYER met5 ;
        RECT -9.180 1200.340 1208.860 1203.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1205.860 -3.820 1208.860 1203.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 21.520 -3.820 23.520 1203.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 86.520 -3.820 88.520 99.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 86.520 501.440 88.520 549.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 86.520 951.440 88.520 1203.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 151.520 -3.820 153.520 89.380 ;
    END
    PORT
      LAYER met4 ;
        RECT 151.520 513.180 153.520 539.380 ;
    END
    PORT
      LAYER met4 ;
        RECT 151.520 963.180 153.520 1203.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 216.520 -3.820 218.520 99.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 216.520 501.440 218.520 549.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 216.520 951.440 218.520 1203.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 281.520 -3.820 283.520 99.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 281.520 501.440 283.520 549.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 281.520 951.440 283.520 1136.855 ;
    END
    PORT
      LAYER met4 ;
        RECT 281.520 1159.415 283.520 1203.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 346.520 -3.820 348.520 99.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 346.520 501.440 348.520 549.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 346.520 951.440 348.520 1203.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 411.520 -3.820 413.520 99.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 411.520 501.440 413.520 549.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 411.520 951.440 413.520 1203.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 476.520 -3.820 478.520 99.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 476.520 501.440 478.520 549.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 476.520 951.440 478.520 1203.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 541.520 -3.820 543.520 1203.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 606.520 -3.820 608.520 1203.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 671.520 -3.820 673.520 1203.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 736.520 -3.820 738.520 1203.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 801.520 -3.820 803.520 1203.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 866.520 -3.820 868.520 1203.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 931.520 -3.820 933.520 1203.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 996.520 -3.820 998.520 1203.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1061.520 -3.820 1063.520 1203.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1126.520 -3.820 1128.520 1203.340 ;
    END
    PORT
      LAYER met4 ;
        RECT 1191.520 -3.820 1193.520 1203.340 ;
    END
    PORT
      LAYER met5 ;
        RECT -9.180 26.880 1208.860 28.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -9.180 91.880 1208.860 93.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -9.180 156.880 166.200 158.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -9.180 221.880 66.420 223.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -9.180 286.880 66.420 288.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -9.180 351.880 66.420 353.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -9.180 416.880 66.420 418.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -9.180 481.880 1208.860 483.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -9.180 546.880 66.420 548.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -9.180 611.880 166.200 613.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -9.180 676.880 166.200 678.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -9.180 741.880 166.200 743.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -9.180 806.880 66.420 808.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -9.180 871.880 66.420 873.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -9.180 936.880 66.420 938.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -9.180 1001.880 1208.860 1003.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -9.180 1066.880 1208.860 1068.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -9.180 1131.880 1208.860 1133.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 353.160 676.880 1208.860 678.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 353.160 741.880 1208.860 743.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 506.200 156.880 1208.860 158.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 506.200 611.880 1208.860 613.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 526.320 221.880 1208.860 223.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 526.320 286.880 1208.860 288.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 526.320 351.880 1208.860 353.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 526.320 416.880 1208.860 418.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 526.320 546.880 1208.860 548.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 526.320 806.880 1208.860 808.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 526.320 871.880 1208.860 873.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 526.320 936.880 1208.860 938.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 21.520 524.300 543.520 526.300 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 20.330 0.000 20.610 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 31.370 0.000 31.650 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 42.410 0.000 42.690 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 53.450 0.000 53.730 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 163.850 0.000 164.130 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 174.890 0.000 175.170 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 185.930 0.000 186.210 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 196.970 0.000 197.250 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 208.010 0.000 208.290 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 219.050 0.000 219.330 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 230.090 0.000 230.370 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 241.130 0.000 241.410 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 252.170 0.000 252.450 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 263.210 0.000 263.490 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 274.250 0.000 274.530 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 285.290 0.000 285.570 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 296.330 0.000 296.610 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 307.370 0.000 307.650 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 318.410 0.000 318.690 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 329.450 0.000 329.730 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 340.490 0.000 340.770 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 351.530 0.000 351.810 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 362.570 0.000 362.850 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 373.610 0.000 373.890 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 75.530 0.000 75.810 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 384.650 0.000 384.930 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 395.690 0.000 395.970 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 86.570 0.000 86.850 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 97.610 0.000 97.890 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 108.650 0.000 108.930 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 119.690 0.000 119.970 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 130.730 0.000 131.010 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 141.770 0.000 142.050 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 152.810 0.000 153.090 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 406.730 0.000 407.010 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 417.770 0.000 418.050 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.170 0.000 528.450 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 539.210 0.000 539.490 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 550.250 0.000 550.530 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 561.290 0.000 561.570 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 572.330 0.000 572.610 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 583.370 0.000 583.650 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 594.410 0.000 594.690 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.450 0.000 605.730 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 616.490 0.000 616.770 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.530 0.000 627.810 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 428.810 0.000 429.090 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 638.570 0.000 638.850 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 649.610 0.000 649.890 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 660.650 0.000 660.930 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 671.690 0.000 671.970 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 682.730 0.000 683.010 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 693.770 0.000 694.050 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 704.810 0.000 705.090 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 715.850 0.000 716.130 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 726.890 0.000 727.170 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.930 0.000 738.210 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 439.850 0.000 440.130 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 748.970 0.000 749.250 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.010 0.000 760.290 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 450.890 0.000 451.170 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.930 0.000 462.210 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.970 0.000 473.250 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.010 0.000 484.290 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.050 0.000 495.330 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 506.090 0.000 506.370 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 517.130 0.000 517.410 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 771.050 0.000 771.330 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 881.450 0.000 881.730 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 892.490 0.000 892.770 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 903.530 0.000 903.810 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 914.570 0.000 914.850 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 925.610 0.000 925.890 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 936.650 0.000 936.930 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 947.690 0.000 947.970 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 958.730 0.000 959.010 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 969.770 0.000 970.050 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 980.810 0.000 981.090 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.090 0.000 782.370 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 991.850 0.000 992.130 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1002.890 0.000 1003.170 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1013.930 0.000 1014.210 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1024.970 0.000 1025.250 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1036.010 0.000 1036.290 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1047.050 0.000 1047.330 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1058.090 0.000 1058.370 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1069.130 0.000 1069.410 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1080.170 0.000 1080.450 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1091.210 0.000 1091.490 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 793.130 0.000 793.410 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1102.250 0.000 1102.530 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1113.290 0.000 1113.570 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 804.170 0.000 804.450 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 815.210 0.000 815.490 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 826.250 0.000 826.530 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 837.290 0.000 837.570 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 848.330 0.000 848.610 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 859.370 0.000 859.650 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 870.410 0.000 870.690 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1124.330 0.000 1124.610 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1135.370 0.000 1135.650 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1146.410 0.000 1146.690 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1157.450 0.000 1157.730 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1168.490 0.000 1168.770 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1179.530 0.000 1179.810 4.000 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1194.160 1188.725 ;
      LAYER met1 ;
        RECT 4.520 9.220 1194.550 1188.880 ;
      LAYER met2 ;
        RECT 4.580 4.280 1194.530 1188.825 ;
        RECT 4.580 4.000 20.050 4.280 ;
        RECT 20.890 4.000 31.090 4.280 ;
        RECT 31.930 4.000 42.130 4.280 ;
        RECT 42.970 4.000 53.170 4.280 ;
        RECT 54.010 4.000 64.210 4.280 ;
        RECT 65.050 4.000 75.250 4.280 ;
        RECT 76.090 4.000 86.290 4.280 ;
        RECT 87.130 4.000 97.330 4.280 ;
        RECT 98.170 4.000 108.370 4.280 ;
        RECT 109.210 4.000 119.410 4.280 ;
        RECT 120.250 4.000 130.450 4.280 ;
        RECT 131.290 4.000 141.490 4.280 ;
        RECT 142.330 4.000 152.530 4.280 ;
        RECT 153.370 4.000 163.570 4.280 ;
        RECT 164.410 4.000 174.610 4.280 ;
        RECT 175.450 4.000 185.650 4.280 ;
        RECT 186.490 4.000 196.690 4.280 ;
        RECT 197.530 4.000 207.730 4.280 ;
        RECT 208.570 4.000 218.770 4.280 ;
        RECT 219.610 4.000 229.810 4.280 ;
        RECT 230.650 4.000 240.850 4.280 ;
        RECT 241.690 4.000 251.890 4.280 ;
        RECT 252.730 4.000 262.930 4.280 ;
        RECT 263.770 4.000 273.970 4.280 ;
        RECT 274.810 4.000 285.010 4.280 ;
        RECT 285.850 4.000 296.050 4.280 ;
        RECT 296.890 4.000 307.090 4.280 ;
        RECT 307.930 4.000 318.130 4.280 ;
        RECT 318.970 4.000 329.170 4.280 ;
        RECT 330.010 4.000 340.210 4.280 ;
        RECT 341.050 4.000 351.250 4.280 ;
        RECT 352.090 4.000 362.290 4.280 ;
        RECT 363.130 4.000 373.330 4.280 ;
        RECT 374.170 4.000 384.370 4.280 ;
        RECT 385.210 4.000 395.410 4.280 ;
        RECT 396.250 4.000 406.450 4.280 ;
        RECT 407.290 4.000 417.490 4.280 ;
        RECT 418.330 4.000 428.530 4.280 ;
        RECT 429.370 4.000 439.570 4.280 ;
        RECT 440.410 4.000 450.610 4.280 ;
        RECT 451.450 4.000 461.650 4.280 ;
        RECT 462.490 4.000 472.690 4.280 ;
        RECT 473.530 4.000 483.730 4.280 ;
        RECT 484.570 4.000 494.770 4.280 ;
        RECT 495.610 4.000 505.810 4.280 ;
        RECT 506.650 4.000 516.850 4.280 ;
        RECT 517.690 4.000 527.890 4.280 ;
        RECT 528.730 4.000 538.930 4.280 ;
        RECT 539.770 4.000 549.970 4.280 ;
        RECT 550.810 4.000 561.010 4.280 ;
        RECT 561.850 4.000 572.050 4.280 ;
        RECT 572.890 4.000 583.090 4.280 ;
        RECT 583.930 4.000 594.130 4.280 ;
        RECT 594.970 4.000 605.170 4.280 ;
        RECT 606.010 4.000 616.210 4.280 ;
        RECT 617.050 4.000 627.250 4.280 ;
        RECT 628.090 4.000 638.290 4.280 ;
        RECT 639.130 4.000 649.330 4.280 ;
        RECT 650.170 4.000 660.370 4.280 ;
        RECT 661.210 4.000 671.410 4.280 ;
        RECT 672.250 4.000 682.450 4.280 ;
        RECT 683.290 4.000 693.490 4.280 ;
        RECT 694.330 4.000 704.530 4.280 ;
        RECT 705.370 4.000 715.570 4.280 ;
        RECT 716.410 4.000 726.610 4.280 ;
        RECT 727.450 4.000 737.650 4.280 ;
        RECT 738.490 4.000 748.690 4.280 ;
        RECT 749.530 4.000 759.730 4.280 ;
        RECT 760.570 4.000 770.770 4.280 ;
        RECT 771.610 4.000 781.810 4.280 ;
        RECT 782.650 4.000 792.850 4.280 ;
        RECT 793.690 4.000 803.890 4.280 ;
        RECT 804.730 4.000 814.930 4.280 ;
        RECT 815.770 4.000 825.970 4.280 ;
        RECT 826.810 4.000 837.010 4.280 ;
        RECT 837.850 4.000 848.050 4.280 ;
        RECT 848.890 4.000 859.090 4.280 ;
        RECT 859.930 4.000 870.130 4.280 ;
        RECT 870.970 4.000 881.170 4.280 ;
        RECT 882.010 4.000 892.210 4.280 ;
        RECT 893.050 4.000 903.250 4.280 ;
        RECT 904.090 4.000 914.290 4.280 ;
        RECT 915.130 4.000 925.330 4.280 ;
        RECT 926.170 4.000 936.370 4.280 ;
        RECT 937.210 4.000 947.410 4.280 ;
        RECT 948.250 4.000 958.450 4.280 ;
        RECT 959.290 4.000 969.490 4.280 ;
        RECT 970.330 4.000 980.530 4.280 ;
        RECT 981.370 4.000 991.570 4.280 ;
        RECT 992.410 4.000 1002.610 4.280 ;
        RECT 1003.450 4.000 1013.650 4.280 ;
        RECT 1014.490 4.000 1024.690 4.280 ;
        RECT 1025.530 4.000 1035.730 4.280 ;
        RECT 1036.570 4.000 1046.770 4.280 ;
        RECT 1047.610 4.000 1057.810 4.280 ;
        RECT 1058.650 4.000 1068.850 4.280 ;
        RECT 1069.690 4.000 1079.890 4.280 ;
        RECT 1080.730 4.000 1090.930 4.280 ;
        RECT 1091.770 4.000 1101.970 4.280 ;
        RECT 1102.810 4.000 1113.010 4.280 ;
        RECT 1113.850 4.000 1124.050 4.280 ;
        RECT 1124.890 4.000 1135.090 4.280 ;
        RECT 1135.930 4.000 1146.130 4.280 ;
        RECT 1146.970 4.000 1157.170 4.280 ;
        RECT 1158.010 4.000 1168.210 4.280 ;
        RECT 1169.050 4.000 1179.250 4.280 ;
        RECT 1180.090 4.000 1194.530 4.280 ;
      LAYER met3 ;
        RECT 2.150 1167.920 1196.000 1188.805 ;
        RECT 4.400 1166.520 1196.000 1167.920 ;
        RECT 2.150 1165.200 1196.000 1166.520 ;
        RECT 2.150 1163.800 1195.600 1165.200 ;
        RECT 2.150 1143.440 1196.000 1163.800 ;
        RECT 2.150 1142.040 1195.600 1143.440 ;
        RECT 2.150 1138.000 1196.000 1142.040 ;
        RECT 4.400 1136.600 1196.000 1138.000 ;
        RECT 2.150 1121.680 1196.000 1136.600 ;
        RECT 2.150 1120.280 1195.600 1121.680 ;
        RECT 2.150 1108.080 1196.000 1120.280 ;
        RECT 4.400 1106.680 1196.000 1108.080 ;
        RECT 2.150 1099.920 1196.000 1106.680 ;
        RECT 2.150 1098.520 1195.600 1099.920 ;
        RECT 2.150 1078.160 1196.000 1098.520 ;
        RECT 4.400 1076.760 1195.600 1078.160 ;
        RECT 2.150 1056.400 1196.000 1076.760 ;
        RECT 2.150 1055.000 1195.600 1056.400 ;
        RECT 2.150 1048.240 1196.000 1055.000 ;
        RECT 4.400 1046.840 1196.000 1048.240 ;
        RECT 2.150 1034.640 1196.000 1046.840 ;
        RECT 2.150 1033.240 1195.600 1034.640 ;
        RECT 2.150 1018.320 1196.000 1033.240 ;
        RECT 4.400 1016.920 1196.000 1018.320 ;
        RECT 2.150 1012.880 1196.000 1016.920 ;
        RECT 2.150 1011.480 1195.600 1012.880 ;
        RECT 2.150 991.120 1196.000 1011.480 ;
        RECT 2.150 989.720 1195.600 991.120 ;
        RECT 2.150 988.400 1196.000 989.720 ;
        RECT 4.400 987.000 1196.000 988.400 ;
        RECT 2.150 969.360 1196.000 987.000 ;
        RECT 2.150 967.960 1195.600 969.360 ;
        RECT 2.150 958.480 1196.000 967.960 ;
        RECT 4.400 957.080 1196.000 958.480 ;
        RECT 2.150 947.600 1196.000 957.080 ;
        RECT 2.150 946.200 1195.600 947.600 ;
        RECT 2.150 928.560 1196.000 946.200 ;
        RECT 4.400 927.160 1196.000 928.560 ;
        RECT 2.150 925.840 1196.000 927.160 ;
        RECT 2.150 924.440 1195.600 925.840 ;
        RECT 2.150 904.080 1196.000 924.440 ;
        RECT 2.150 902.680 1195.600 904.080 ;
        RECT 2.150 898.640 1196.000 902.680 ;
        RECT 4.400 897.240 1196.000 898.640 ;
        RECT 2.150 882.320 1196.000 897.240 ;
        RECT 2.150 880.920 1195.600 882.320 ;
        RECT 2.150 868.720 1196.000 880.920 ;
        RECT 4.400 867.320 1196.000 868.720 ;
        RECT 2.150 860.560 1196.000 867.320 ;
        RECT 2.150 859.160 1195.600 860.560 ;
        RECT 2.150 838.800 1196.000 859.160 ;
        RECT 4.400 837.400 1195.600 838.800 ;
        RECT 2.150 817.040 1196.000 837.400 ;
        RECT 2.150 815.640 1195.600 817.040 ;
        RECT 2.150 808.880 1196.000 815.640 ;
        RECT 4.400 807.480 1196.000 808.880 ;
        RECT 2.150 795.280 1196.000 807.480 ;
        RECT 2.150 793.880 1195.600 795.280 ;
        RECT 2.150 778.960 1196.000 793.880 ;
        RECT 4.400 777.560 1196.000 778.960 ;
        RECT 2.150 773.520 1196.000 777.560 ;
        RECT 2.150 772.120 1195.600 773.520 ;
        RECT 2.150 751.760 1196.000 772.120 ;
        RECT 2.150 750.360 1195.600 751.760 ;
        RECT 2.150 749.040 1196.000 750.360 ;
        RECT 4.400 747.640 1196.000 749.040 ;
        RECT 2.150 730.000 1196.000 747.640 ;
        RECT 2.150 728.600 1195.600 730.000 ;
        RECT 2.150 719.120 1196.000 728.600 ;
        RECT 4.400 717.720 1196.000 719.120 ;
        RECT 2.150 708.240 1196.000 717.720 ;
        RECT 2.150 706.840 1195.600 708.240 ;
        RECT 2.150 689.200 1196.000 706.840 ;
        RECT 4.400 687.800 1196.000 689.200 ;
        RECT 2.150 686.480 1196.000 687.800 ;
        RECT 2.150 685.080 1195.600 686.480 ;
        RECT 2.150 664.720 1196.000 685.080 ;
        RECT 2.150 663.320 1195.600 664.720 ;
        RECT 2.150 659.280 1196.000 663.320 ;
        RECT 4.400 657.880 1196.000 659.280 ;
        RECT 2.150 642.960 1196.000 657.880 ;
        RECT 2.150 641.560 1195.600 642.960 ;
        RECT 2.150 629.360 1196.000 641.560 ;
        RECT 4.400 627.960 1196.000 629.360 ;
        RECT 2.150 621.200 1196.000 627.960 ;
        RECT 2.150 619.800 1195.600 621.200 ;
        RECT 2.150 599.440 1196.000 619.800 ;
        RECT 4.400 598.040 1195.600 599.440 ;
        RECT 2.150 577.680 1196.000 598.040 ;
        RECT 2.150 576.280 1195.600 577.680 ;
        RECT 2.150 569.520 1196.000 576.280 ;
        RECT 4.400 568.120 1196.000 569.520 ;
        RECT 2.150 555.920 1196.000 568.120 ;
        RECT 2.150 554.520 1195.600 555.920 ;
        RECT 2.150 539.600 1196.000 554.520 ;
        RECT 4.400 538.200 1196.000 539.600 ;
        RECT 2.150 534.160 1196.000 538.200 ;
        RECT 2.150 532.760 1195.600 534.160 ;
        RECT 2.150 512.400 1196.000 532.760 ;
        RECT 2.150 511.000 1195.600 512.400 ;
        RECT 2.150 509.680 1196.000 511.000 ;
        RECT 4.400 508.280 1196.000 509.680 ;
        RECT 2.150 490.640 1196.000 508.280 ;
        RECT 2.150 489.240 1195.600 490.640 ;
        RECT 2.150 479.760 1196.000 489.240 ;
        RECT 4.400 478.360 1196.000 479.760 ;
        RECT 2.150 468.880 1196.000 478.360 ;
        RECT 2.150 467.480 1195.600 468.880 ;
        RECT 2.150 449.840 1196.000 467.480 ;
        RECT 4.400 448.440 1196.000 449.840 ;
        RECT 2.150 447.120 1196.000 448.440 ;
        RECT 2.150 445.720 1195.600 447.120 ;
        RECT 2.150 425.360 1196.000 445.720 ;
        RECT 2.150 423.960 1195.600 425.360 ;
        RECT 2.150 419.920 1196.000 423.960 ;
        RECT 4.400 418.520 1196.000 419.920 ;
        RECT 2.150 403.600 1196.000 418.520 ;
        RECT 2.150 402.200 1195.600 403.600 ;
        RECT 2.150 390.000 1196.000 402.200 ;
        RECT 4.400 388.600 1196.000 390.000 ;
        RECT 2.150 381.840 1196.000 388.600 ;
        RECT 2.150 380.440 1195.600 381.840 ;
        RECT 2.150 360.080 1196.000 380.440 ;
        RECT 4.400 358.680 1195.600 360.080 ;
        RECT 2.150 338.320 1196.000 358.680 ;
        RECT 2.150 336.920 1195.600 338.320 ;
        RECT 2.150 330.160 1196.000 336.920 ;
        RECT 4.400 328.760 1196.000 330.160 ;
        RECT 2.150 316.560 1196.000 328.760 ;
        RECT 2.150 315.160 1195.600 316.560 ;
        RECT 2.150 300.240 1196.000 315.160 ;
        RECT 4.400 298.840 1196.000 300.240 ;
        RECT 2.150 294.800 1196.000 298.840 ;
        RECT 2.150 293.400 1195.600 294.800 ;
        RECT 2.150 273.040 1196.000 293.400 ;
        RECT 2.150 271.640 1195.600 273.040 ;
        RECT 2.150 270.320 1196.000 271.640 ;
        RECT 4.400 268.920 1196.000 270.320 ;
        RECT 2.150 251.280 1196.000 268.920 ;
        RECT 2.150 249.880 1195.600 251.280 ;
        RECT 2.150 240.400 1196.000 249.880 ;
        RECT 4.400 239.000 1196.000 240.400 ;
        RECT 2.150 229.520 1196.000 239.000 ;
        RECT 2.150 228.120 1195.600 229.520 ;
        RECT 2.150 210.480 1196.000 228.120 ;
        RECT 4.400 209.080 1196.000 210.480 ;
        RECT 2.150 207.760 1196.000 209.080 ;
        RECT 2.150 206.360 1195.600 207.760 ;
        RECT 2.150 186.000 1196.000 206.360 ;
        RECT 2.150 184.600 1195.600 186.000 ;
        RECT 2.150 180.560 1196.000 184.600 ;
        RECT 4.400 179.160 1196.000 180.560 ;
        RECT 2.150 164.240 1196.000 179.160 ;
        RECT 2.150 162.840 1195.600 164.240 ;
        RECT 2.150 150.640 1196.000 162.840 ;
        RECT 4.400 149.240 1196.000 150.640 ;
        RECT 2.150 142.480 1196.000 149.240 ;
        RECT 2.150 141.080 1195.600 142.480 ;
        RECT 2.150 120.720 1196.000 141.080 ;
        RECT 4.400 119.320 1195.600 120.720 ;
        RECT 2.150 98.960 1196.000 119.320 ;
        RECT 2.150 97.560 1195.600 98.960 ;
        RECT 2.150 90.800 1196.000 97.560 ;
        RECT 4.400 89.400 1196.000 90.800 ;
        RECT 2.150 77.200 1196.000 89.400 ;
        RECT 2.150 75.800 1195.600 77.200 ;
        RECT 2.150 60.880 1196.000 75.800 ;
        RECT 4.400 59.480 1196.000 60.880 ;
        RECT 2.150 55.440 1196.000 59.480 ;
        RECT 2.150 54.040 1195.600 55.440 ;
        RECT 2.150 33.680 1196.000 54.040 ;
        RECT 2.150 32.280 1195.600 33.680 ;
        RECT 2.150 30.960 1196.000 32.280 ;
        RECT 4.400 29.560 1196.000 30.960 ;
        RECT 2.150 10.715 1196.000 29.560 ;
      LAYER met4 ;
        RECT 53.655 99.980 69.120 1152.890 ;
        RECT 71.920 951.040 86.120 1152.890 ;
        RECT 88.920 1141.205 151.120 1152.890 ;
        RECT 88.920 951.040 134.120 1141.205 ;
        RECT 136.920 962.780 151.120 1141.205 ;
        RECT 153.920 962.780 199.120 1152.890 ;
        RECT 136.920 951.040 199.120 962.780 ;
        RECT 201.920 951.040 216.120 1152.890 ;
        RECT 218.920 951.040 264.120 1152.890 ;
        RECT 266.920 1137.255 329.120 1152.890 ;
        RECT 266.920 951.040 281.120 1137.255 ;
        RECT 283.920 951.040 329.120 1137.255 ;
        RECT 331.920 951.040 346.120 1152.890 ;
        RECT 348.920 951.040 394.120 1152.890 ;
        RECT 396.920 951.040 411.120 1152.890 ;
        RECT 413.920 1137.255 476.120 1152.890 ;
        RECT 413.920 951.040 459.120 1137.255 ;
        RECT 461.920 951.040 476.120 1137.255 ;
        RECT 478.920 951.040 524.120 1152.890 ;
        RECT 71.920 549.800 524.120 951.040 ;
        RECT 71.920 501.040 86.120 549.800 ;
        RECT 88.920 501.040 134.120 549.800 ;
        RECT 136.920 539.780 199.120 549.800 ;
        RECT 136.920 512.780 151.120 539.780 ;
        RECT 153.920 512.780 199.120 539.780 ;
        RECT 136.920 501.040 199.120 512.780 ;
        RECT 201.920 501.040 216.120 549.800 ;
        RECT 218.920 501.040 264.120 549.800 ;
        RECT 266.920 501.040 281.120 549.800 ;
        RECT 283.920 501.040 329.120 549.800 ;
        RECT 331.920 501.040 346.120 549.800 ;
        RECT 348.920 501.040 394.120 549.800 ;
        RECT 396.920 501.040 411.120 549.800 ;
        RECT 413.920 501.040 459.120 549.800 ;
        RECT 461.920 501.040 476.120 549.800 ;
        RECT 478.920 501.040 524.120 549.800 ;
        RECT 71.920 99.980 524.120 501.040 ;
        RECT 526.920 99.980 541.120 1152.890 ;
        RECT 543.920 99.980 589.120 1152.890 ;
        RECT 591.920 99.980 606.120 1152.890 ;
        RECT 608.920 99.980 627.490 1152.890 ;
      LAYER met5 ;
        RECT 79.620 1135.480 627.500 1152.900 ;
        RECT 79.620 1118.480 627.500 1130.280 ;
        RECT 79.620 1070.480 627.500 1113.280 ;
        RECT 79.620 1053.480 627.500 1065.280 ;
        RECT 79.620 1005.480 627.500 1048.280 ;
        RECT 79.620 988.480 627.500 1000.280 ;
        RECT 79.620 940.480 627.500 983.280 ;
        RECT 79.620 935.280 524.720 940.480 ;
        RECT 79.620 923.480 627.500 935.280 ;
        RECT 79.620 918.280 524.720 923.480 ;
        RECT 79.620 875.480 627.500 918.280 ;
        RECT 79.620 870.280 524.720 875.480 ;
        RECT 79.620 858.480 627.500 870.280 ;
        RECT 79.620 853.280 522.920 858.480 ;
        RECT 79.620 810.480 627.500 853.280 ;
        RECT 79.620 805.280 524.720 810.480 ;
        RECT 79.620 793.480 627.500 805.280 ;
        RECT 167.800 788.280 351.560 793.480 ;
        RECT 79.620 745.480 627.500 788.280 ;
        RECT 167.800 740.280 351.560 745.480 ;
        RECT 79.620 728.480 627.500 740.280 ;
        RECT 167.800 723.280 351.560 728.480 ;
        RECT 79.620 680.480 627.500 723.280 ;
        RECT 167.800 675.280 351.560 680.480 ;
        RECT 79.620 663.480 627.500 675.280 ;
        RECT 79.620 658.280 522.920 663.480 ;
        RECT 79.620 615.480 627.500 658.280 ;
        RECT 167.800 610.280 504.600 615.480 ;
        RECT 79.620 598.480 627.500 610.280 ;
        RECT 79.620 593.280 524.720 598.480 ;
        RECT 79.620 550.480 627.500 593.280 ;
        RECT 79.620 545.280 524.720 550.480 ;
        RECT 79.620 533.480 627.500 545.280 ;
        RECT 79.620 527.900 627.500 528.280 ;
        RECT 545.120 522.700 627.500 527.900 ;
        RECT 79.620 485.480 627.500 522.700 ;
        RECT 79.620 468.480 627.500 480.280 ;
        RECT 79.620 463.280 524.720 468.480 ;
        RECT 79.620 420.480 627.500 463.280 ;
        RECT 79.620 415.280 524.720 420.480 ;
        RECT 79.620 403.480 627.500 415.280 ;
        RECT 79.620 398.280 524.720 403.480 ;
        RECT 79.620 355.480 627.500 398.280 ;
        RECT 79.620 350.280 524.720 355.480 ;
        RECT 79.620 338.480 627.500 350.280 ;
        RECT 79.620 333.280 524.720 338.480 ;
        RECT 79.620 290.480 627.500 333.280 ;
        RECT 79.620 285.280 524.720 290.480 ;
        RECT 79.620 273.480 627.500 285.280 ;
        RECT 167.800 268.280 351.560 273.480 ;
        RECT 79.620 225.480 627.500 268.280 ;
        RECT 79.620 220.280 524.720 225.480 ;
        RECT 79.620 208.480 627.500 220.280 ;
        RECT 167.800 203.280 394.930 208.480 ;
        RECT 79.620 160.480 627.500 203.280 ;
        RECT 167.800 155.280 504.600 160.480 ;
        RECT 79.620 143.480 627.500 155.280 ;
        RECT 79.620 138.280 522.920 143.480 ;
        RECT 79.620 99.980 627.500 138.280 ;
  END
END signal_generator
END LIBRARY

