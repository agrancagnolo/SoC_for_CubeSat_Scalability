VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wb_buttons_leds
  CLASS BLOCK ;
  FOREIGN wb_buttons_leds ;
  ORIGIN 0.000 0.000 ;
  SIZE 2800.000 BY 500.000 ;
  PIN buttons[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 20.440 2800.000 21.040 ;
    END
  END buttons[0]
  PIN buttons[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 58.520 2800.000 59.120 ;
    END
  END buttons[1]
  PIN buttons[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 96.600 2800.000 97.200 ;
    END
  END buttons[2]
  PIN led_enb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 172.760 2800.000 173.360 ;
    END
  END led_enb[0]
  PIN led_enb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 248.920 2800.000 249.520 ;
    END
  END led_enb[1]
  PIN led_enb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 325.080 2800.000 325.680 ;
    END
  END led_enb[2]
  PIN led_enb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 401.240 2800.000 401.840 ;
    END
  END led_enb[3]
  PIN led_enb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 477.400 2800.000 478.000 ;
    END
  END led_enb[4]
  PIN led_enb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.040 4.000 374.640 ;
    END
  END led_enb[5]
  PIN led_enb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 208.120 4.000 208.720 ;
    END
  END led_enb[6]
  PIN led_enb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.200 4.000 42.800 ;
    END
  END led_enb[7]
  PIN leds[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 134.680 2800.000 135.280 ;
    END
  END leds[0]
  PIN leds[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 210.840 2800.000 211.440 ;
    END
  END leds[1]
  PIN leds[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 287.000 2800.000 287.600 ;
    END
  END leds[2]
  PIN leds[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 363.160 2800.000 363.760 ;
    END
  END leds[3]
  PIN leds[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 439.320 2800.000 439.920 ;
    END
  END leds[4]
  PIN leds[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 457.000 4.000 457.600 ;
    END
  END leds[5]
  PIN leds[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 291.080 4.000 291.680 ;
    END
  END leds[6]
  PIN leds[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.160 4.000 125.760 ;
    END
  END leds[7]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 1557.040 10.640 1558.640 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 1710.640 10.640 1712.240 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 1864.240 10.640 1865.840 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 2017.840 10.640 2019.440 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 2171.440 10.640 2173.040 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 2325.040 10.640 2326.640 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 2478.640 10.640 2480.240 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 2632.240 10.640 2633.840 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 2785.840 10.640 2787.440 487.120 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 1633.840 10.640 1635.440 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 1787.440 10.640 1789.040 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 1941.040 10.640 1942.640 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 2094.640 10.640 2096.240 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 2248.240 10.640 2249.840 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 2401.840 10.640 2403.440 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 2555.440 10.640 2557.040 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 2709.040 10.640 2710.640 487.120 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 56.210 0.000 56.490 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 83.350 0.000 83.630 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 191.910 0.000 192.190 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1006.110 0.000 1006.390 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1087.530 0.000 1087.810 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1168.950 0.000 1169.230 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1250.370 0.000 1250.650 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1331.790 0.000 1332.070 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1413.210 0.000 1413.490 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1494.630 0.000 1494.910 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1576.050 0.000 1576.330 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1657.470 0.000 1657.750 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1738.890 0.000 1739.170 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 273.330 0.000 273.610 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1820.310 0.000 1820.590 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1901.730 0.000 1902.010 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1983.150 0.000 1983.430 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 2064.570 0.000 2064.850 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 2145.990 0.000 2146.270 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 2227.410 0.000 2227.690 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 2308.830 0.000 2309.110 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 2390.250 0.000 2390.530 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 2471.670 0.000 2471.950 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 2553.090 0.000 2553.370 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 354.750 0.000 355.030 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 2634.510 0.000 2634.790 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 2715.930 0.000 2716.210 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 436.170 0.000 436.450 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 517.590 0.000 517.870 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 599.010 0.000 599.290 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 680.430 0.000 680.710 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 761.850 0.000 762.130 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 843.270 0.000 843.550 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 924.690 0.000 924.970 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 110.490 0.000 110.770 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 219.050 0.000 219.330 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1033.250 0.000 1033.530 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1114.670 0.000 1114.950 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1196.090 0.000 1196.370 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1277.510 0.000 1277.790 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1358.930 0.000 1359.210 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1440.350 0.000 1440.630 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1521.770 0.000 1522.050 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1603.190 0.000 1603.470 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1684.610 0.000 1684.890 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1766.030 0.000 1766.310 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 300.470 0.000 300.750 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1847.450 0.000 1847.730 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1928.870 0.000 1929.150 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2010.290 0.000 2010.570 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2091.710 0.000 2091.990 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2173.130 0.000 2173.410 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2254.550 0.000 2254.830 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2335.970 0.000 2336.250 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2417.390 0.000 2417.670 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2498.810 0.000 2499.090 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2580.230 0.000 2580.510 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 381.890 0.000 382.170 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2661.650 0.000 2661.930 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2743.070 0.000 2743.350 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 463.310 0.000 463.590 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 544.730 0.000 545.010 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 626.150 0.000 626.430 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 707.570 0.000 707.850 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 788.990 0.000 789.270 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 870.410 0.000 870.690 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 951.830 0.000 952.110 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 246.190 0.000 246.470 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1060.390 0.000 1060.670 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1141.810 0.000 1142.090 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1223.230 0.000 1223.510 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1304.650 0.000 1304.930 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1386.070 0.000 1386.350 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1467.490 0.000 1467.770 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1548.910 0.000 1549.190 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1630.330 0.000 1630.610 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1711.750 0.000 1712.030 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1793.170 0.000 1793.450 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 327.610 0.000 327.890 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1874.590 0.000 1874.870 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1956.010 0.000 1956.290 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2037.430 0.000 2037.710 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2118.850 0.000 2119.130 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2200.270 0.000 2200.550 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2281.690 0.000 2281.970 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2363.110 0.000 2363.390 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2444.530 0.000 2444.810 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2525.950 0.000 2526.230 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2607.370 0.000 2607.650 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 409.030 0.000 409.310 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2688.790 0.000 2689.070 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2770.210 0.000 2770.490 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 490.450 0.000 490.730 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 571.870 0.000 572.150 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 653.290 0.000 653.570 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 734.710 0.000 734.990 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 816.130 0.000 816.410 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 897.550 0.000 897.830 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 978.970 0.000 979.250 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 137.630 0.000 137.910 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 164.770 0.000 165.050 4.000 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 2794.040 486.965 ;
      LAYER met1 ;
        RECT 4.670 6.840 2794.040 487.120 ;
      LAYER met2 ;
        RECT 4.690 4.280 2792.570 487.065 ;
        RECT 4.690 3.670 28.790 4.280 ;
        RECT 29.630 3.670 55.930 4.280 ;
        RECT 56.770 3.670 83.070 4.280 ;
        RECT 83.910 3.670 110.210 4.280 ;
        RECT 111.050 3.670 137.350 4.280 ;
        RECT 138.190 3.670 164.490 4.280 ;
        RECT 165.330 3.670 191.630 4.280 ;
        RECT 192.470 3.670 218.770 4.280 ;
        RECT 219.610 3.670 245.910 4.280 ;
        RECT 246.750 3.670 273.050 4.280 ;
        RECT 273.890 3.670 300.190 4.280 ;
        RECT 301.030 3.670 327.330 4.280 ;
        RECT 328.170 3.670 354.470 4.280 ;
        RECT 355.310 3.670 381.610 4.280 ;
        RECT 382.450 3.670 408.750 4.280 ;
        RECT 409.590 3.670 435.890 4.280 ;
        RECT 436.730 3.670 463.030 4.280 ;
        RECT 463.870 3.670 490.170 4.280 ;
        RECT 491.010 3.670 517.310 4.280 ;
        RECT 518.150 3.670 544.450 4.280 ;
        RECT 545.290 3.670 571.590 4.280 ;
        RECT 572.430 3.670 598.730 4.280 ;
        RECT 599.570 3.670 625.870 4.280 ;
        RECT 626.710 3.670 653.010 4.280 ;
        RECT 653.850 3.670 680.150 4.280 ;
        RECT 680.990 3.670 707.290 4.280 ;
        RECT 708.130 3.670 734.430 4.280 ;
        RECT 735.270 3.670 761.570 4.280 ;
        RECT 762.410 3.670 788.710 4.280 ;
        RECT 789.550 3.670 815.850 4.280 ;
        RECT 816.690 3.670 842.990 4.280 ;
        RECT 843.830 3.670 870.130 4.280 ;
        RECT 870.970 3.670 897.270 4.280 ;
        RECT 898.110 3.670 924.410 4.280 ;
        RECT 925.250 3.670 951.550 4.280 ;
        RECT 952.390 3.670 978.690 4.280 ;
        RECT 979.530 3.670 1005.830 4.280 ;
        RECT 1006.670 3.670 1032.970 4.280 ;
        RECT 1033.810 3.670 1060.110 4.280 ;
        RECT 1060.950 3.670 1087.250 4.280 ;
        RECT 1088.090 3.670 1114.390 4.280 ;
        RECT 1115.230 3.670 1141.530 4.280 ;
        RECT 1142.370 3.670 1168.670 4.280 ;
        RECT 1169.510 3.670 1195.810 4.280 ;
        RECT 1196.650 3.670 1222.950 4.280 ;
        RECT 1223.790 3.670 1250.090 4.280 ;
        RECT 1250.930 3.670 1277.230 4.280 ;
        RECT 1278.070 3.670 1304.370 4.280 ;
        RECT 1305.210 3.670 1331.510 4.280 ;
        RECT 1332.350 3.670 1358.650 4.280 ;
        RECT 1359.490 3.670 1385.790 4.280 ;
        RECT 1386.630 3.670 1412.930 4.280 ;
        RECT 1413.770 3.670 1440.070 4.280 ;
        RECT 1440.910 3.670 1467.210 4.280 ;
        RECT 1468.050 3.670 1494.350 4.280 ;
        RECT 1495.190 3.670 1521.490 4.280 ;
        RECT 1522.330 3.670 1548.630 4.280 ;
        RECT 1549.470 3.670 1575.770 4.280 ;
        RECT 1576.610 3.670 1602.910 4.280 ;
        RECT 1603.750 3.670 1630.050 4.280 ;
        RECT 1630.890 3.670 1657.190 4.280 ;
        RECT 1658.030 3.670 1684.330 4.280 ;
        RECT 1685.170 3.670 1711.470 4.280 ;
        RECT 1712.310 3.670 1738.610 4.280 ;
        RECT 1739.450 3.670 1765.750 4.280 ;
        RECT 1766.590 3.670 1792.890 4.280 ;
        RECT 1793.730 3.670 1820.030 4.280 ;
        RECT 1820.870 3.670 1847.170 4.280 ;
        RECT 1848.010 3.670 1874.310 4.280 ;
        RECT 1875.150 3.670 1901.450 4.280 ;
        RECT 1902.290 3.670 1928.590 4.280 ;
        RECT 1929.430 3.670 1955.730 4.280 ;
        RECT 1956.570 3.670 1982.870 4.280 ;
        RECT 1983.710 3.670 2010.010 4.280 ;
        RECT 2010.850 3.670 2037.150 4.280 ;
        RECT 2037.990 3.670 2064.290 4.280 ;
        RECT 2065.130 3.670 2091.430 4.280 ;
        RECT 2092.270 3.670 2118.570 4.280 ;
        RECT 2119.410 3.670 2145.710 4.280 ;
        RECT 2146.550 3.670 2172.850 4.280 ;
        RECT 2173.690 3.670 2199.990 4.280 ;
        RECT 2200.830 3.670 2227.130 4.280 ;
        RECT 2227.970 3.670 2254.270 4.280 ;
        RECT 2255.110 3.670 2281.410 4.280 ;
        RECT 2282.250 3.670 2308.550 4.280 ;
        RECT 2309.390 3.670 2335.690 4.280 ;
        RECT 2336.530 3.670 2362.830 4.280 ;
        RECT 2363.670 3.670 2389.970 4.280 ;
        RECT 2390.810 3.670 2417.110 4.280 ;
        RECT 2417.950 3.670 2444.250 4.280 ;
        RECT 2445.090 3.670 2471.390 4.280 ;
        RECT 2472.230 3.670 2498.530 4.280 ;
        RECT 2499.370 3.670 2525.670 4.280 ;
        RECT 2526.510 3.670 2552.810 4.280 ;
        RECT 2553.650 3.670 2579.950 4.280 ;
        RECT 2580.790 3.670 2607.090 4.280 ;
        RECT 2607.930 3.670 2634.230 4.280 ;
        RECT 2635.070 3.670 2661.370 4.280 ;
        RECT 2662.210 3.670 2688.510 4.280 ;
        RECT 2689.350 3.670 2715.650 4.280 ;
        RECT 2716.490 3.670 2742.790 4.280 ;
        RECT 2743.630 3.670 2769.930 4.280 ;
        RECT 2770.770 3.670 2792.570 4.280 ;
      LAYER met3 ;
        RECT 4.000 478.400 2796.000 487.045 ;
        RECT 4.000 477.000 2795.600 478.400 ;
        RECT 4.000 458.000 2796.000 477.000 ;
        RECT 4.400 456.600 2796.000 458.000 ;
        RECT 4.000 440.320 2796.000 456.600 ;
        RECT 4.000 438.920 2795.600 440.320 ;
        RECT 4.000 402.240 2796.000 438.920 ;
        RECT 4.000 400.840 2795.600 402.240 ;
        RECT 4.000 375.040 2796.000 400.840 ;
        RECT 4.400 373.640 2796.000 375.040 ;
        RECT 4.000 364.160 2796.000 373.640 ;
        RECT 4.000 362.760 2795.600 364.160 ;
        RECT 4.000 326.080 2796.000 362.760 ;
        RECT 4.000 324.680 2795.600 326.080 ;
        RECT 4.000 292.080 2796.000 324.680 ;
        RECT 4.400 290.680 2796.000 292.080 ;
        RECT 4.000 288.000 2796.000 290.680 ;
        RECT 4.000 286.600 2795.600 288.000 ;
        RECT 4.000 249.920 2796.000 286.600 ;
        RECT 4.000 248.520 2795.600 249.920 ;
        RECT 4.000 211.840 2796.000 248.520 ;
        RECT 4.000 210.440 2795.600 211.840 ;
        RECT 4.000 209.120 2796.000 210.440 ;
        RECT 4.400 207.720 2796.000 209.120 ;
        RECT 4.000 173.760 2796.000 207.720 ;
        RECT 4.000 172.360 2795.600 173.760 ;
        RECT 4.000 135.680 2796.000 172.360 ;
        RECT 4.000 134.280 2795.600 135.680 ;
        RECT 4.000 126.160 2796.000 134.280 ;
        RECT 4.400 124.760 2796.000 126.160 ;
        RECT 4.000 97.600 2796.000 124.760 ;
        RECT 4.000 96.200 2795.600 97.600 ;
        RECT 4.000 59.520 2796.000 96.200 ;
        RECT 4.000 58.120 2795.600 59.520 ;
        RECT 4.000 43.200 2796.000 58.120 ;
        RECT 4.400 41.800 2796.000 43.200 ;
        RECT 4.000 21.440 2796.000 41.800 ;
        RECT 4.000 20.040 2795.600 21.440 ;
        RECT 4.000 10.715 2796.000 20.040 ;
  END
END wb_buttons_leds
END LIBRARY

