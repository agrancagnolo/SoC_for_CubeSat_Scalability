* NGSPICE file created from Mixer.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_01v8_Y6SADL a_n210_n1149# a_n50_n1063# a_50_n975# a_n108_n975#
X0 a_50_n975# a_n50_n1063# a_n108_n975# a_n210_n1149# sky130_fd_pr__nfet_01v8 ad=2.8275 pd=20.08 as=2.8275 ps=20.08 w=9.75 l=0.5
.ends

.subckt sky130_fd_pr__nfet_01v8_Y6FLEL a_n210_n1149# a_n50_n1063# a_50_n975# a_n108_n975#
X0 a_50_n975# a_n50_n1063# a_n108_n975# a_n210_n1149# sky130_fd_pr__nfet_01v8 ad=2.8275 pd=20.08 as=2.8275 ps=20.08 w=9.75 l=0.5
.ends

.subckt sky130_fd_pr__nfet_01v8_PZKCVB a_n50_n1038# a_50_n950# a_n108_n950# a_n210_n1124#
X0 a_50_n950# a_n50_n1038# a_n108_n950# a_n210_n1124# sky130_fd_pr__nfet_01v8 ad=2.755 pd=19.58 as=2.755 ps=19.58 w=9.5 l=0.5
.ends

.subckt sky130_fd_pr__nfet_01v8_PMG9RB a_n50_n1038# a_50_n950# a_n108_n950# a_n210_n1124#
X0 a_50_n950# a_n50_n1038# a_n108_n950# a_n210_n1124# sky130_fd_pr__nfet_01v8 ad=2.755 pd=19.58 as=2.755 ps=19.58 w=9.5 l=0.5
.ends

.subckt sky130_fd_pr__nfet_01v8_8XPPYK a_n123_n1515# a_n65_n1570# a_65_n1515# a_n225_n1689#
X0 a_65_n1515# a_n65_n1570# a_n123_n1515# a_n225_n1689# sky130_fd_pr__nfet_01v8 ad=4.3935 pd=30.88 as=4.3935 ps=30.88 w=15.15 l=0.65
.ends

.subckt sky130_fd_pr__nfet_01v8_Z6VF7Q a_n50_n1038# a_50_n950# a_n108_n950# a_n210_n1124#
X0 a_50_n950# a_n50_n1038# a_n108_n950# a_n210_n1124# sky130_fd_pr__nfet_01v8 ad=2.755 pd=19.58 as=2.755 ps=19.58 w=9.5 l=0.5
.ends

.subckt sky130_fd_pr__nfet_01v8_Z9V85Y a_n50_n1038# a_50_n950# a_n108_n950# a_n210_n1124#
X0 a_50_n950# a_n50_n1038# a_n108_n950# a_n210_n1124# sky130_fd_pr__nfet_01v8 ad=2.755 pd=19.58 as=2.755 ps=19.58 w=9.5 l=0.5
.ends

.subckt sky130_fd_pr__nfet_01v8_VJM6P6 a_n210_n1149# a_n50_n1063# a_50_n975# a_n108_n975#
X0 a_50_n975# a_n50_n1063# a_n108_n975# a_n210_n1149# sky130_fd_pr__nfet_01v8 ad=2.8275 pd=20.08 as=2.8275 ps=20.08 w=9.75 l=0.5
.ends

.subckt sky130_fd_pr__nfet_01v8_HQ3Y9H a_n210_n1149# a_n50_n1063# a_50_n975# a_n108_n975#
X0 a_50_n975# a_n50_n1063# a_n108_n975# a_n210_n1149# sky130_fd_pr__nfet_01v8 ad=2.8275 pd=20.08 as=2.8275 ps=20.08 w=9.75 l=0.5
.ends

.subckt sky130_fd_pr__pfet_01v8_JCZH34 a_n50_n967# a_n108_n870# w_n246_n1089# a_50_n870#
X0 a_50_n870# a_n50_n967# a_n108_n870# w_n246_n1089# sky130_fd_pr__pfet_01v8 ad=2.523 pd=17.98 as=2.523 ps=17.98 w=8.7 l=0.5
.ends

.subckt sky130_fd_pr__pfet_01v8_9F3ELE a_n50_n297# a_50_n200# a_n108_n200# w_n246_n419#
X0 a_50_n200# a_n50_n297# a_n108_n200# w_n246_n419# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
.ends

.subckt sky130_fd_pr__pfet_01v8_4F365H a_n50_n297# a_50_n200# a_n108_n200# w_n246_n419#
X0 a_50_n200# a_n50_n297# a_n108_n200# w_n246_n419# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
.ends

.subckt sky130_fd_pr__pfet_01v8_53Y4NB a_n50_n967# a_n108_n870# w_n246_n1089# a_50_n870#
X0 a_50_n870# a_n50_n967# a_n108_n870# w_n246_n1089# sky130_fd_pr__pfet_01v8 ad=2.523 pd=17.98 as=2.523 ps=17.98 w=8.7 l=0.5
.ends

.subckt Mixer vdd gnd vlo- out- vlo+ vbias2 vbias3 vrf+ vrf- vtail vbias1 out+
XXM1 gnd vrf+ m1_5180_850# m1_4048_1162# sky130_fd_pr__nfet_01v8_Y6SADL
XXM2 gnd vrf- m1_5180_850# m1_4436_2196# sky130_fd_pr__nfet_01v8_Y6FLEL
XXM3 vlo- m1_962_656# out+ gnd sky130_fd_pr__nfet_01v8_PZKCVB
XXM4 vlo+ m1_962_656# out- gnd sky130_fd_pr__nfet_01v8_PMG9RB
XXMTAIL m1_5180_850# vtail gnd gnd sky130_fd_pr__nfet_01v8_8XPPYK
XXM5 vlo+ m1_2744_894# out+ gnd sky130_fd_pr__nfet_01v8_Z6VF7Q
XXM6 vlo- m1_2744_894# out- gnd sky130_fd_pr__nfet_01v8_Z9V85Y
XXM7 gnd vbias1 m1_4048_1162# m1_962_656# sky130_fd_pr__nfet_01v8_VJM6P6
XXM8 gnd vbias1 m1_4436_2196# m1_2744_894# sky130_fd_pr__nfet_01v8_HQ3Y9H
XXM9 vbias2 out+ vdd vdd sky130_fd_pr__pfet_01v8_JCZH34
XXMci2 vbias3 vdd m1_2744_894# vdd sky130_fd_pr__pfet_01v8_9F3ELE
XXMci1 vbias3 vdd m1_962_656# vdd sky130_fd_pr__pfet_01v8_4F365H
XXM10 vbias2 out- vdd vdd sky130_fd_pr__pfet_01v8_53Y4NB
.ends

