VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO signal_generator
  CLASS BLOCK ;
  FOREIGN signal_generator ;
  ORIGIN 0.000 0.000 ;
  SIZE 1200.000 BY 1200.000 ;
  PIN io_analog[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 32.680 1200.000 33.280 ;
    END
  END io_analog[0]
  PIN io_analog[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 250.280 1200.000 250.880 ;
    END
  END io_analog[10]
  PIN io_analog[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 54.440 1200.000 55.040 ;
    END
  END io_analog[1]
  PIN io_analog[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 76.200 1200.000 76.800 ;
    END
  END io_analog[2]
  PIN io_analog[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 97.960 1200.000 98.560 ;
    END
  END io_analog[3]
  PIN io_analog[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 119.720 1200.000 120.320 ;
    END
  END io_analog[4]
  PIN io_analog[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 141.480 1200.000 142.080 ;
    END
  END io_analog[5]
  PIN io_analog[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1196.000 163.240 1200.000 163.840 ;
    END
  END io_analog[6]
  PIN io_analog[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 1196.000 185.000 1200.000 185.600 ;
    END
  END io_analog[7]
  PIN io_analog[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1196.000 206.760 1200.000 207.360 ;
    END
  END io_analog[8]
  PIN io_analog[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1196.000 228.520 1200.000 229.120 ;
    END
  END io_analog[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 272.040 1200.000 272.640 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 924.840 1200.000 925.440 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 990.120 1200.000 990.720 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1055.400 1200.000 1056.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1120.680 1200.000 1121.280 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1166.920 4.000 1167.520 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1077.160 4.000 1077.760 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 987.400 4.000 988.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 897.640 4.000 898.240 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 807.880 4.000 808.480 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 718.120 4.000 718.720 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 337.320 1200.000 337.920 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 628.360 4.000 628.960 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 538.600 4.000 539.200 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 448.840 4.000 449.440 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 359.080 4.000 359.680 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 269.320 4.000 269.920 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 179.560 4.000 180.160 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.800 4.000 90.400 ;
    END
  END io_in[26]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 402.600 1200.000 403.200 ;
    END
  END io_in[2]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 467.880 1200.000 468.480 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 533.160 1200.000 533.760 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 598.440 1200.000 599.040 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 663.720 1200.000 664.320 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 729.000 1200.000 729.600 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 794.280 1200.000 794.880 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 859.560 1200.000 860.160 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 315.560 1200.000 316.160 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 968.360 1200.000 968.960 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1033.640 1200.000 1034.240 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1098.920 1200.000 1099.520 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1164.200 1200.000 1164.800 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1107.080 4.000 1107.680 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1017.320 4.000 1017.920 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 927.560 4.000 928.160 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 837.800 4.000 838.400 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 748.040 4.000 748.640 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 658.280 4.000 658.880 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 380.840 1200.000 381.440 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 568.520 4.000 569.120 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 478.760 4.000 479.360 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 389.000 4.000 389.600 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.240 4.000 299.840 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 209.480 4.000 210.080 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.720 4.000 120.320 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.960 4.000 30.560 ;
    END
  END io_oeb[26]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 446.120 1200.000 446.720 ;
    END
  END io_oeb[2]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 511.400 1200.000 512.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 576.680 1200.000 577.280 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 641.960 1200.000 642.560 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 707.240 1200.000 707.840 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 772.520 1200.000 773.120 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 837.800 1200.000 838.400 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 903.080 1200.000 903.680 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 293.800 1200.000 294.400 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 1196.000 946.600 1200.000 947.200 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1011.880 1200.000 1012.480 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1077.160 1200.000 1077.760 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1142.440 1200.000 1143.040 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1137.000 4.000 1137.600 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1047.240 4.000 1047.840 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 957.480 4.000 958.080 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 867.720 4.000 868.320 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 777.960 4.000 778.560 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 688.200 4.000 688.800 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 359.080 1200.000 359.680 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 598.440 4.000 599.040 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 508.680 4.000 509.280 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 418.920 4.000 419.520 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 329.160 4.000 329.760 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 239.400 4.000 240.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.880 4.000 60.480 ;
    END
  END io_out[26]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 424.360 1200.000 424.960 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 489.640 1200.000 490.240 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 554.920 1200.000 555.520 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 620.200 1200.000 620.800 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 685.480 1200.000 686.080 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 1196.000 750.760 1200.000 751.360 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 1196.000 816.040 1200.000 816.640 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 1196.000 881.320 1200.000 881.920 ;
    END
  END io_out[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.120 0.880 3.120 1187.760 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.120 0.880 1189.900 3.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.120 1184.760 1189.900 1187.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 1186.900 0.880 1189.900 1187.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 9.120 -3.820 11.120 1192.460 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.120 -3.820 76.120 1192.460 ;
    END
    PORT
      LAYER met4 ;
        RECT 139.120 -3.820 141.120 1192.460 ;
    END
    PORT
      LAYER met4 ;
        RECT 204.120 -3.820 206.120 99.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 204.120 501.440 206.120 549.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 204.120 951.440 206.120 1192.460 ;
    END
    PORT
      LAYER met4 ;
        RECT 269.120 -3.820 271.120 99.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 269.120 501.440 271.120 549.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 269.120 951.440 271.120 1192.460 ;
    END
    PORT
      LAYER met4 ;
        RECT 334.120 -3.820 336.120 99.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 334.120 501.440 336.120 549.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 334.120 951.440 336.120 1192.460 ;
    END
    PORT
      LAYER met4 ;
        RECT 399.120 -3.820 401.120 99.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 399.120 501.440 401.120 549.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 399.120 951.440 401.120 1192.460 ;
    END
    PORT
      LAYER met4 ;
        RECT 464.120 -3.820 466.120 99.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 464.120 501.440 466.120 549.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 464.120 951.440 466.120 1192.460 ;
    END
    PORT
      LAYER met4 ;
        RECT 529.120 -3.820 531.120 99.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 529.120 501.440 531.120 549.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 529.120 951.440 531.120 1192.460 ;
    END
    PORT
      LAYER met4 ;
        RECT 594.120 -3.820 596.120 1192.460 ;
    END
    PORT
      LAYER met4 ;
        RECT 659.120 -3.820 661.120 1192.460 ;
    END
    PORT
      LAYER met4 ;
        RECT 724.120 -3.820 726.120 1192.460 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.120 -3.820 791.120 1192.460 ;
    END
    PORT
      LAYER met4 ;
        RECT 854.120 -3.820 856.120 1192.460 ;
    END
    PORT
      LAYER met4 ;
        RECT 919.120 -3.820 921.120 1192.460 ;
    END
    PORT
      LAYER met4 ;
        RECT 984.120 -3.820 986.120 1192.460 ;
    END
    PORT
      LAYER met4 ;
        RECT 1049.120 -3.820 1051.120 680.805 ;
    END
    PORT
      LAYER met4 ;
        RECT 1049.120 703.365 1051.120 1078.805 ;
    END
    PORT
      LAYER met4 ;
        RECT 1049.120 1101.360 1051.120 1192.460 ;
    END
    PORT
      LAYER met4 ;
        RECT 1114.120 -3.820 1116.120 1192.460 ;
    END
    PORT
      LAYER met5 ;
        RECT -4.580 9.880 1194.600 11.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -4.580 74.880 1194.600 76.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -4.580 139.880 136.420 141.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -4.580 204.880 236.200 206.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -4.580 269.880 236.200 271.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -4.580 334.880 136.420 336.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -4.580 399.880 136.420 401.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -4.580 464.880 136.420 466.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -4.580 529.880 1194.600 531.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -4.580 594.880 136.420 596.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -4.580 659.880 136.420 661.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -4.580 724.880 236.200 726.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -4.580 789.880 236.200 791.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -4.580 854.880 136.420 856.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -4.580 919.880 136.420 921.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -4.580 984.880 1194.600 986.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -4.580 1049.880 1194.600 1051.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -4.580 1114.880 1194.600 1116.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 423.160 269.880 1194.600 271.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 423.160 724.880 1194.600 726.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 423.160 789.880 1194.600 791.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 466.530 204.880 1194.600 206.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 596.320 139.880 1194.600 141.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 596.320 334.880 1194.600 336.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 596.320 399.880 1194.600 401.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 596.320 464.880 1194.600 466.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 596.320 594.880 1194.600 596.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 596.320 659.880 1194.600 661.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 596.320 854.880 1194.600 856.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 596.320 919.880 1194.600 921.880 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -4.580 -3.820 -1.580 1192.460 ;
    END
    PORT
      LAYER met5 ;
        RECT -4.580 -3.820 1194.600 -0.820 ;
    END
    PORT
      LAYER met5 ;
        RECT -4.580 1189.460 1194.600 1192.460 ;
    END
    PORT
      LAYER met4 ;
        RECT 1191.600 -3.820 1194.600 1192.460 ;
    END
    PORT
      LAYER met4 ;
        RECT 26.120 -3.820 28.120 1192.460 ;
    END
    PORT
      LAYER met4 ;
        RECT 91.120 -3.820 93.120 1192.460 ;
    END
    PORT
      LAYER met4 ;
        RECT 156.120 -3.820 158.120 99.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 156.120 501.440 158.120 549.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 156.120 951.440 158.120 1192.460 ;
    END
    PORT
      LAYER met4 ;
        RECT 221.120 -3.820 223.120 89.380 ;
    END
    PORT
      LAYER met4 ;
        RECT 221.120 513.180 223.120 539.380 ;
    END
    PORT
      LAYER met4 ;
        RECT 221.120 963.180 223.120 1192.460 ;
    END
    PORT
      LAYER met4 ;
        RECT 286.120 -3.820 288.120 99.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 286.120 501.440 288.120 549.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 286.120 951.440 288.120 1192.460 ;
    END
    PORT
      LAYER met4 ;
        RECT 351.120 -3.820 353.120 99.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 351.120 501.440 353.120 549.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 351.120 951.440 353.120 1192.460 ;
    END
    PORT
      LAYER met4 ;
        RECT 416.120 -3.820 418.120 99.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 416.120 501.440 418.120 549.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 416.120 951.440 418.120 1192.460 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.120 -3.820 483.120 99.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.120 501.440 483.120 549.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.120 951.440 483.120 1192.460 ;
    END
    PORT
      LAYER met4 ;
        RECT 546.120 -3.820 548.120 99.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 546.120 501.440 548.120 549.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 546.120 951.440 548.120 1192.460 ;
    END
    PORT
      LAYER met4 ;
        RECT 611.120 -3.820 613.120 1192.460 ;
    END
    PORT
      LAYER met4 ;
        RECT 676.120 -3.820 678.120 1192.460 ;
    END
    PORT
      LAYER met4 ;
        RECT 741.120 -3.820 743.120 1192.460 ;
    END
    PORT
      LAYER met4 ;
        RECT 806.120 -3.820 808.120 1192.460 ;
    END
    PORT
      LAYER met4 ;
        RECT 871.120 -3.820 873.120 1192.460 ;
    END
    PORT
      LAYER met4 ;
        RECT 936.120 -3.820 938.120 1192.460 ;
    END
    PORT
      LAYER met4 ;
        RECT 1001.120 -3.820 1003.120 1192.460 ;
    END
    PORT
      LAYER met4 ;
        RECT 1066.120 -3.820 1068.120 1192.460 ;
    END
    PORT
      LAYER met4 ;
        RECT 1131.120 -3.820 1133.120 1192.460 ;
    END
    PORT
      LAYER met5 ;
        RECT -4.580 26.880 1194.600 28.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -4.580 91.880 1194.600 93.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -4.580 156.880 236.200 158.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -4.580 221.880 136.420 223.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -4.580 286.880 136.420 288.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -4.580 351.880 136.420 353.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -4.580 416.880 136.420 418.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -4.580 481.880 1194.600 483.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -4.580 546.880 136.420 548.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -4.580 611.880 236.200 613.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -4.580 676.880 236.200 678.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -4.580 741.880 236.200 743.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -4.580 806.880 136.420 808.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -4.580 871.880 136.420 873.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -4.580 936.880 136.420 938.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -4.580 1001.880 1194.600 1003.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -4.580 1066.880 1194.600 1068.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -4.580 1131.880 1194.600 1133.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 423.160 676.880 1194.600 678.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 423.160 741.880 1194.600 743.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 576.200 156.880 1194.600 158.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 576.200 611.880 1194.600 613.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 596.320 221.880 1194.600 223.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 596.320 286.880 1194.600 288.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 596.320 351.880 1194.600 353.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 596.320 416.880 1194.600 418.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 596.320 546.880 1194.600 548.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 596.320 806.880 1194.600 808.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 596.320 871.880 1194.600 873.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 596.320 936.880 1194.600 938.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 91.120 524.300 613.120 526.300 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 20.330 0.000 20.610 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 31.370 0.000 31.650 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 42.410 0.000 42.690 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 53.450 0.000 53.730 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 163.850 0.000 164.130 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 174.890 0.000 175.170 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 185.930 0.000 186.210 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 196.970 0.000 197.250 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 208.010 0.000 208.290 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 219.050 0.000 219.330 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 230.090 0.000 230.370 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 241.130 0.000 241.410 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 252.170 0.000 252.450 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 263.210 0.000 263.490 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 274.250 0.000 274.530 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 285.290 0.000 285.570 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 296.330 0.000 296.610 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 307.370 0.000 307.650 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 318.410 0.000 318.690 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 329.450 0.000 329.730 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 340.490 0.000 340.770 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 351.530 0.000 351.810 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 362.570 0.000 362.850 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 373.610 0.000 373.890 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 75.530 0.000 75.810 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 384.650 0.000 384.930 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 395.690 0.000 395.970 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 86.570 0.000 86.850 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 97.610 0.000 97.890 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 108.650 0.000 108.930 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 119.690 0.000 119.970 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 130.730 0.000 131.010 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 141.770 0.000 142.050 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 152.810 0.000 153.090 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 406.730 0.000 407.010 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 417.770 0.000 418.050 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.170 0.000 528.450 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 539.210 0.000 539.490 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 550.250 0.000 550.530 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 561.290 0.000 561.570 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 572.330 0.000 572.610 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 583.370 0.000 583.650 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 594.410 0.000 594.690 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.450 0.000 605.730 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 616.490 0.000 616.770 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.530 0.000 627.810 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 428.810 0.000 429.090 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 638.570 0.000 638.850 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 649.610 0.000 649.890 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 660.650 0.000 660.930 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 671.690 0.000 671.970 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 682.730 0.000 683.010 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 693.770 0.000 694.050 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 704.810 0.000 705.090 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 715.850 0.000 716.130 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 726.890 0.000 727.170 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.930 0.000 738.210 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 439.850 0.000 440.130 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 748.970 0.000 749.250 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.010 0.000 760.290 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 450.890 0.000 451.170 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.930 0.000 462.210 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.970 0.000 473.250 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.010 0.000 484.290 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.050 0.000 495.330 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 506.090 0.000 506.370 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 517.130 0.000 517.410 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 771.050 0.000 771.330 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 881.450 0.000 881.730 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 892.490 0.000 892.770 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 903.530 0.000 903.810 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 914.570 0.000 914.850 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 925.610 0.000 925.890 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 936.650 0.000 936.930 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 947.690 0.000 947.970 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 958.730 0.000 959.010 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 969.770 0.000 970.050 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 980.810 0.000 981.090 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.090 0.000 782.370 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 991.850 0.000 992.130 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1002.890 0.000 1003.170 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1013.930 0.000 1014.210 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1024.970 0.000 1025.250 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1036.010 0.000 1036.290 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1047.050 0.000 1047.330 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1058.090 0.000 1058.370 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1069.130 0.000 1069.410 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1080.170 0.000 1080.450 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1091.210 0.000 1091.490 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 793.130 0.000 793.410 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1102.250 0.000 1102.530 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1113.290 0.000 1113.570 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 804.170 0.000 804.450 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 815.210 0.000 815.490 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 826.250 0.000 826.530 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 837.290 0.000 837.570 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 848.330 0.000 848.610 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 859.370 0.000 859.650 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 870.410 0.000 870.690 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1124.330 0.000 1124.610 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1135.370 0.000 1135.650 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1146.410 0.000 1146.690 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1157.450 0.000 1157.730 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1168.490 0.000 1168.770 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1179.530 0.000 1179.810 4.000 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 10.120 10.795 1179.900 1177.845 ;
      LAYER met1 ;
        RECT 6.510 9.220 1187.650 1178.000 ;
      LAYER met2 ;
        RECT 6.530 4.280 1187.630 1177.945 ;
        RECT 6.530 3.670 20.050 4.280 ;
        RECT 20.890 3.670 31.090 4.280 ;
        RECT 31.930 3.670 42.130 4.280 ;
        RECT 42.970 3.670 53.170 4.280 ;
        RECT 54.010 3.670 64.210 4.280 ;
        RECT 65.050 3.670 75.250 4.280 ;
        RECT 76.090 3.670 86.290 4.280 ;
        RECT 87.130 3.670 97.330 4.280 ;
        RECT 98.170 3.670 108.370 4.280 ;
        RECT 109.210 3.670 119.410 4.280 ;
        RECT 120.250 3.670 130.450 4.280 ;
        RECT 131.290 3.670 141.490 4.280 ;
        RECT 142.330 3.670 152.530 4.280 ;
        RECT 153.370 3.670 163.570 4.280 ;
        RECT 164.410 3.670 174.610 4.280 ;
        RECT 175.450 3.670 185.650 4.280 ;
        RECT 186.490 3.670 196.690 4.280 ;
        RECT 197.530 3.670 207.730 4.280 ;
        RECT 208.570 3.670 218.770 4.280 ;
        RECT 219.610 3.670 229.810 4.280 ;
        RECT 230.650 3.670 240.850 4.280 ;
        RECT 241.690 3.670 251.890 4.280 ;
        RECT 252.730 3.670 262.930 4.280 ;
        RECT 263.770 3.670 273.970 4.280 ;
        RECT 274.810 3.670 285.010 4.280 ;
        RECT 285.850 3.670 296.050 4.280 ;
        RECT 296.890 3.670 307.090 4.280 ;
        RECT 307.930 3.670 318.130 4.280 ;
        RECT 318.970 3.670 329.170 4.280 ;
        RECT 330.010 3.670 340.210 4.280 ;
        RECT 341.050 3.670 351.250 4.280 ;
        RECT 352.090 3.670 362.290 4.280 ;
        RECT 363.130 3.670 373.330 4.280 ;
        RECT 374.170 3.670 384.370 4.280 ;
        RECT 385.210 3.670 395.410 4.280 ;
        RECT 396.250 3.670 406.450 4.280 ;
        RECT 407.290 3.670 417.490 4.280 ;
        RECT 418.330 3.670 428.530 4.280 ;
        RECT 429.370 3.670 439.570 4.280 ;
        RECT 440.410 3.670 450.610 4.280 ;
        RECT 451.450 3.670 461.650 4.280 ;
        RECT 462.490 3.670 472.690 4.280 ;
        RECT 473.530 3.670 483.730 4.280 ;
        RECT 484.570 3.670 494.770 4.280 ;
        RECT 495.610 3.670 505.810 4.280 ;
        RECT 506.650 3.670 516.850 4.280 ;
        RECT 517.690 3.670 527.890 4.280 ;
        RECT 528.730 3.670 538.930 4.280 ;
        RECT 539.770 3.670 549.970 4.280 ;
        RECT 550.810 3.670 561.010 4.280 ;
        RECT 561.850 3.670 572.050 4.280 ;
        RECT 572.890 3.670 583.090 4.280 ;
        RECT 583.930 3.670 594.130 4.280 ;
        RECT 594.970 3.670 605.170 4.280 ;
        RECT 606.010 3.670 616.210 4.280 ;
        RECT 617.050 3.670 627.250 4.280 ;
        RECT 628.090 3.670 638.290 4.280 ;
        RECT 639.130 3.670 649.330 4.280 ;
        RECT 650.170 3.670 660.370 4.280 ;
        RECT 661.210 3.670 671.410 4.280 ;
        RECT 672.250 3.670 682.450 4.280 ;
        RECT 683.290 3.670 693.490 4.280 ;
        RECT 694.330 3.670 704.530 4.280 ;
        RECT 705.370 3.670 715.570 4.280 ;
        RECT 716.410 3.670 726.610 4.280 ;
        RECT 727.450 3.670 737.650 4.280 ;
        RECT 738.490 3.670 748.690 4.280 ;
        RECT 749.530 3.670 759.730 4.280 ;
        RECT 760.570 3.670 770.770 4.280 ;
        RECT 771.610 3.670 781.810 4.280 ;
        RECT 782.650 3.670 792.850 4.280 ;
        RECT 793.690 3.670 803.890 4.280 ;
        RECT 804.730 3.670 814.930 4.280 ;
        RECT 815.770 3.670 825.970 4.280 ;
        RECT 826.810 3.670 837.010 4.280 ;
        RECT 837.850 3.670 848.050 4.280 ;
        RECT 848.890 3.670 859.090 4.280 ;
        RECT 859.930 3.670 870.130 4.280 ;
        RECT 870.970 3.670 881.170 4.280 ;
        RECT 882.010 3.670 892.210 4.280 ;
        RECT 893.050 3.670 903.250 4.280 ;
        RECT 904.090 3.670 914.290 4.280 ;
        RECT 915.130 3.670 925.330 4.280 ;
        RECT 926.170 3.670 936.370 4.280 ;
        RECT 937.210 3.670 947.410 4.280 ;
        RECT 948.250 3.670 958.450 4.280 ;
        RECT 959.290 3.670 969.490 4.280 ;
        RECT 970.330 3.670 980.530 4.280 ;
        RECT 981.370 3.670 991.570 4.280 ;
        RECT 992.410 3.670 1002.610 4.280 ;
        RECT 1003.450 3.670 1013.650 4.280 ;
        RECT 1014.490 3.670 1024.690 4.280 ;
        RECT 1025.530 3.670 1035.730 4.280 ;
        RECT 1036.570 3.670 1046.770 4.280 ;
        RECT 1047.610 3.670 1057.810 4.280 ;
        RECT 1058.650 3.670 1068.850 4.280 ;
        RECT 1069.690 3.670 1079.890 4.280 ;
        RECT 1080.730 3.670 1090.930 4.280 ;
        RECT 1091.770 3.670 1101.970 4.280 ;
        RECT 1102.810 3.670 1113.010 4.280 ;
        RECT 1113.850 3.670 1124.050 4.280 ;
        RECT 1124.890 3.670 1135.090 4.280 ;
        RECT 1135.930 3.670 1146.130 4.280 ;
        RECT 1146.970 3.670 1157.170 4.280 ;
        RECT 1158.010 3.670 1168.210 4.280 ;
        RECT 1169.050 3.670 1179.250 4.280 ;
        RECT 1180.090 3.670 1187.630 4.280 ;
      LAYER met3 ;
        RECT 4.000 1167.920 1196.000 1177.925 ;
        RECT 4.400 1166.520 1196.000 1167.920 ;
        RECT 4.000 1165.200 1196.000 1166.520 ;
        RECT 4.000 1163.800 1195.600 1165.200 ;
        RECT 4.000 1143.440 1196.000 1163.800 ;
        RECT 4.000 1142.040 1195.600 1143.440 ;
        RECT 4.000 1138.000 1196.000 1142.040 ;
        RECT 4.400 1136.600 1196.000 1138.000 ;
        RECT 4.000 1121.680 1196.000 1136.600 ;
        RECT 4.000 1120.280 1195.600 1121.680 ;
        RECT 4.000 1108.080 1196.000 1120.280 ;
        RECT 4.400 1106.680 1196.000 1108.080 ;
        RECT 4.000 1099.920 1196.000 1106.680 ;
        RECT 4.000 1098.520 1195.600 1099.920 ;
        RECT 4.000 1078.160 1196.000 1098.520 ;
        RECT 4.400 1076.760 1195.600 1078.160 ;
        RECT 4.000 1056.400 1196.000 1076.760 ;
        RECT 4.000 1055.000 1195.600 1056.400 ;
        RECT 4.000 1048.240 1196.000 1055.000 ;
        RECT 4.400 1046.840 1196.000 1048.240 ;
        RECT 4.000 1034.640 1196.000 1046.840 ;
        RECT 4.000 1033.240 1195.600 1034.640 ;
        RECT 4.000 1018.320 1196.000 1033.240 ;
        RECT 4.400 1016.920 1196.000 1018.320 ;
        RECT 4.000 1012.880 1196.000 1016.920 ;
        RECT 4.000 1011.480 1195.600 1012.880 ;
        RECT 4.000 991.120 1196.000 1011.480 ;
        RECT 4.000 989.720 1195.600 991.120 ;
        RECT 4.000 988.400 1196.000 989.720 ;
        RECT 4.400 987.000 1196.000 988.400 ;
        RECT 4.000 969.360 1196.000 987.000 ;
        RECT 4.000 967.960 1195.600 969.360 ;
        RECT 4.000 958.480 1196.000 967.960 ;
        RECT 4.400 957.080 1196.000 958.480 ;
        RECT 4.000 947.600 1196.000 957.080 ;
        RECT 4.000 946.200 1195.600 947.600 ;
        RECT 4.000 928.560 1196.000 946.200 ;
        RECT 4.400 927.160 1196.000 928.560 ;
        RECT 4.000 925.840 1196.000 927.160 ;
        RECT 4.000 924.440 1195.600 925.840 ;
        RECT 4.000 904.080 1196.000 924.440 ;
        RECT 4.000 902.680 1195.600 904.080 ;
        RECT 4.000 898.640 1196.000 902.680 ;
        RECT 4.400 897.240 1196.000 898.640 ;
        RECT 4.000 882.320 1196.000 897.240 ;
        RECT 4.000 880.920 1195.600 882.320 ;
        RECT 4.000 868.720 1196.000 880.920 ;
        RECT 4.400 867.320 1196.000 868.720 ;
        RECT 4.000 860.560 1196.000 867.320 ;
        RECT 4.000 859.160 1195.600 860.560 ;
        RECT 4.000 838.800 1196.000 859.160 ;
        RECT 4.400 837.400 1195.600 838.800 ;
        RECT 4.000 817.040 1196.000 837.400 ;
        RECT 4.000 815.640 1195.600 817.040 ;
        RECT 4.000 808.880 1196.000 815.640 ;
        RECT 4.400 807.480 1196.000 808.880 ;
        RECT 4.000 795.280 1196.000 807.480 ;
        RECT 4.000 793.880 1195.600 795.280 ;
        RECT 4.000 778.960 1196.000 793.880 ;
        RECT 4.400 777.560 1196.000 778.960 ;
        RECT 4.000 773.520 1196.000 777.560 ;
        RECT 4.000 772.120 1195.600 773.520 ;
        RECT 4.000 751.760 1196.000 772.120 ;
        RECT 4.000 750.360 1195.600 751.760 ;
        RECT 4.000 749.040 1196.000 750.360 ;
        RECT 4.400 747.640 1196.000 749.040 ;
        RECT 4.000 730.000 1196.000 747.640 ;
        RECT 4.000 728.600 1195.600 730.000 ;
        RECT 4.000 719.120 1196.000 728.600 ;
        RECT 4.400 717.720 1196.000 719.120 ;
        RECT 4.000 708.240 1196.000 717.720 ;
        RECT 4.000 706.840 1195.600 708.240 ;
        RECT 4.000 689.200 1196.000 706.840 ;
        RECT 4.400 687.800 1196.000 689.200 ;
        RECT 4.000 686.480 1196.000 687.800 ;
        RECT 4.000 685.080 1195.600 686.480 ;
        RECT 4.000 664.720 1196.000 685.080 ;
        RECT 4.000 663.320 1195.600 664.720 ;
        RECT 4.000 659.280 1196.000 663.320 ;
        RECT 4.400 657.880 1196.000 659.280 ;
        RECT 4.000 642.960 1196.000 657.880 ;
        RECT 4.000 641.560 1195.600 642.960 ;
        RECT 4.000 629.360 1196.000 641.560 ;
        RECT 4.400 627.960 1196.000 629.360 ;
        RECT 4.000 621.200 1196.000 627.960 ;
        RECT 4.000 619.800 1195.600 621.200 ;
        RECT 4.000 599.440 1196.000 619.800 ;
        RECT 4.400 598.040 1195.600 599.440 ;
        RECT 4.000 577.680 1196.000 598.040 ;
        RECT 4.000 576.280 1195.600 577.680 ;
        RECT 4.000 569.520 1196.000 576.280 ;
        RECT 4.400 568.120 1196.000 569.520 ;
        RECT 4.000 555.920 1196.000 568.120 ;
        RECT 4.000 554.520 1195.600 555.920 ;
        RECT 4.000 539.600 1196.000 554.520 ;
        RECT 4.400 538.200 1196.000 539.600 ;
        RECT 4.000 534.160 1196.000 538.200 ;
        RECT 4.000 532.760 1195.600 534.160 ;
        RECT 4.000 512.400 1196.000 532.760 ;
        RECT 4.000 511.000 1195.600 512.400 ;
        RECT 4.000 509.680 1196.000 511.000 ;
        RECT 4.400 508.280 1196.000 509.680 ;
        RECT 4.000 490.640 1196.000 508.280 ;
        RECT 4.000 489.240 1195.600 490.640 ;
        RECT 4.000 479.760 1196.000 489.240 ;
        RECT 4.400 478.360 1196.000 479.760 ;
        RECT 4.000 468.880 1196.000 478.360 ;
        RECT 4.000 467.480 1195.600 468.880 ;
        RECT 4.000 449.840 1196.000 467.480 ;
        RECT 4.400 448.440 1196.000 449.840 ;
        RECT 4.000 447.120 1196.000 448.440 ;
        RECT 4.000 445.720 1195.600 447.120 ;
        RECT 4.000 425.360 1196.000 445.720 ;
        RECT 4.000 423.960 1195.600 425.360 ;
        RECT 4.000 419.920 1196.000 423.960 ;
        RECT 4.400 418.520 1196.000 419.920 ;
        RECT 4.000 403.600 1196.000 418.520 ;
        RECT 4.000 402.200 1195.600 403.600 ;
        RECT 4.000 390.000 1196.000 402.200 ;
        RECT 4.400 388.600 1196.000 390.000 ;
        RECT 4.000 381.840 1196.000 388.600 ;
        RECT 4.000 380.440 1195.600 381.840 ;
        RECT 4.000 360.080 1196.000 380.440 ;
        RECT 4.400 358.680 1195.600 360.080 ;
        RECT 4.000 338.320 1196.000 358.680 ;
        RECT 4.000 336.920 1195.600 338.320 ;
        RECT 4.000 330.160 1196.000 336.920 ;
        RECT 4.400 328.760 1196.000 330.160 ;
        RECT 4.000 316.560 1196.000 328.760 ;
        RECT 4.000 315.160 1195.600 316.560 ;
        RECT 4.000 300.240 1196.000 315.160 ;
        RECT 4.400 298.840 1196.000 300.240 ;
        RECT 4.000 294.800 1196.000 298.840 ;
        RECT 4.000 293.400 1195.600 294.800 ;
        RECT 4.000 273.040 1196.000 293.400 ;
        RECT 4.000 271.640 1195.600 273.040 ;
        RECT 4.000 270.320 1196.000 271.640 ;
        RECT 4.400 268.920 1196.000 270.320 ;
        RECT 4.000 251.280 1196.000 268.920 ;
        RECT 4.000 249.880 1195.600 251.280 ;
        RECT 4.000 240.400 1196.000 249.880 ;
        RECT 4.400 239.000 1196.000 240.400 ;
        RECT 4.000 229.520 1196.000 239.000 ;
        RECT 4.000 228.120 1195.600 229.520 ;
        RECT 4.000 210.480 1196.000 228.120 ;
        RECT 4.400 209.080 1196.000 210.480 ;
        RECT 4.000 207.760 1196.000 209.080 ;
        RECT 4.000 206.360 1195.600 207.760 ;
        RECT 4.000 186.000 1196.000 206.360 ;
        RECT 4.000 184.600 1195.600 186.000 ;
        RECT 4.000 180.560 1196.000 184.600 ;
        RECT 4.400 179.160 1196.000 180.560 ;
        RECT 4.000 164.240 1196.000 179.160 ;
        RECT 4.000 162.840 1195.600 164.240 ;
        RECT 4.000 150.640 1196.000 162.840 ;
        RECT 4.400 149.240 1196.000 150.640 ;
        RECT 4.000 142.480 1196.000 149.240 ;
        RECT 4.000 141.080 1195.600 142.480 ;
        RECT 4.000 120.720 1196.000 141.080 ;
        RECT 4.400 119.320 1195.600 120.720 ;
        RECT 4.000 98.960 1196.000 119.320 ;
        RECT 4.000 97.560 1195.600 98.960 ;
        RECT 4.000 90.800 1196.000 97.560 ;
        RECT 4.400 89.400 1196.000 90.800 ;
        RECT 4.000 77.200 1196.000 89.400 ;
        RECT 4.000 75.800 1195.600 77.200 ;
        RECT 4.000 60.880 1196.000 75.800 ;
        RECT 4.400 59.480 1196.000 60.880 ;
        RECT 4.000 55.440 1196.000 59.480 ;
        RECT 4.000 54.040 1195.600 55.440 ;
        RECT 4.000 33.680 1196.000 54.040 ;
        RECT 4.000 32.280 1195.600 33.680 ;
        RECT 4.000 30.960 1196.000 32.280 ;
        RECT 4.400 29.560 1196.000 30.960 ;
        RECT 4.000 10.715 1196.000 29.560 ;
      LAYER met4 ;
        RECT 118.975 83.135 138.720 1090.890 ;
        RECT 141.520 951.040 155.720 1090.890 ;
        RECT 158.520 951.040 203.720 1090.890 ;
        RECT 206.520 962.780 220.720 1090.890 ;
        RECT 223.520 962.780 268.720 1090.890 ;
        RECT 206.520 951.040 268.720 962.780 ;
        RECT 271.520 951.040 285.720 1090.890 ;
        RECT 288.520 951.040 333.720 1090.890 ;
        RECT 336.520 951.040 350.720 1090.890 ;
        RECT 353.520 951.040 398.720 1090.890 ;
        RECT 401.520 951.040 415.720 1090.890 ;
        RECT 418.520 951.040 463.720 1090.890 ;
        RECT 466.520 951.040 480.720 1090.890 ;
        RECT 483.520 951.040 528.720 1090.890 ;
        RECT 531.520 951.040 545.720 1090.890 ;
        RECT 548.520 951.040 593.720 1090.890 ;
        RECT 141.520 549.800 593.720 951.040 ;
        RECT 141.520 501.040 155.720 549.800 ;
        RECT 158.520 501.040 203.720 549.800 ;
        RECT 206.520 539.780 268.720 549.800 ;
        RECT 206.520 512.780 220.720 539.780 ;
        RECT 223.520 512.780 268.720 539.780 ;
        RECT 206.520 501.040 268.720 512.780 ;
        RECT 271.520 501.040 285.720 549.800 ;
        RECT 288.520 501.040 333.720 549.800 ;
        RECT 336.520 501.040 350.720 549.800 ;
        RECT 353.520 501.040 398.720 549.800 ;
        RECT 401.520 501.040 415.720 549.800 ;
        RECT 418.520 501.040 463.720 549.800 ;
        RECT 466.520 501.040 480.720 549.800 ;
        RECT 483.520 501.040 528.720 549.800 ;
        RECT 531.520 501.040 545.720 549.800 ;
        RECT 548.520 501.040 593.720 549.800 ;
        RECT 141.520 99.800 593.720 501.040 ;
        RECT 141.520 83.135 155.720 99.800 ;
        RECT 158.520 83.135 203.720 99.800 ;
        RECT 206.520 89.780 268.720 99.800 ;
        RECT 206.520 83.135 220.720 89.780 ;
        RECT 223.520 83.135 268.720 89.780 ;
        RECT 271.520 83.135 285.720 99.800 ;
        RECT 288.520 83.135 333.720 99.800 ;
        RECT 336.520 83.135 350.720 99.800 ;
        RECT 353.520 83.135 398.720 99.800 ;
        RECT 401.520 83.135 415.720 99.800 ;
        RECT 418.520 83.135 463.720 99.800 ;
        RECT 466.520 83.135 480.720 99.800 ;
        RECT 483.520 83.135 528.720 99.800 ;
        RECT 531.520 83.135 545.720 99.800 ;
        RECT 548.520 83.135 593.720 99.800 ;
        RECT 596.520 83.135 610.720 1090.890 ;
        RECT 613.520 83.135 658.720 1090.890 ;
        RECT 661.520 83.135 675.720 1090.890 ;
        RECT 678.520 83.135 723.720 1090.890 ;
        RECT 726.520 83.135 740.720 1090.890 ;
        RECT 743.520 83.135 788.720 1090.890 ;
        RECT 791.520 83.135 805.720 1090.890 ;
        RECT 808.520 83.135 853.720 1090.890 ;
        RECT 856.520 83.135 870.720 1090.890 ;
        RECT 873.520 83.135 918.720 1090.890 ;
        RECT 921.520 83.135 935.720 1090.890 ;
        RECT 938.520 83.135 983.720 1090.890 ;
        RECT 986.520 83.135 1000.720 1090.890 ;
        RECT 1003.520 1079.205 1065.720 1090.890 ;
        RECT 1003.520 702.965 1048.720 1079.205 ;
        RECT 1051.520 702.965 1065.720 1079.205 ;
        RECT 1003.520 681.205 1065.720 702.965 ;
        RECT 1003.520 83.135 1048.720 681.205 ;
        RECT 1051.520 83.135 1065.720 681.205 ;
        RECT 1068.520 83.135 1092.490 1090.890 ;
      LAYER met5 ;
        RECT 149.620 1070.480 1092.500 1090.900 ;
        RECT 149.620 1053.480 1092.500 1065.280 ;
        RECT 149.620 1005.480 1092.500 1048.280 ;
        RECT 149.620 988.480 1092.500 1000.280 ;
        RECT 149.620 940.480 1092.500 983.280 ;
        RECT 149.620 935.280 594.720 940.480 ;
        RECT 149.620 923.480 1092.500 935.280 ;
        RECT 149.620 918.280 594.720 923.480 ;
        RECT 149.620 875.480 1092.500 918.280 ;
        RECT 149.620 870.280 594.720 875.480 ;
        RECT 149.620 858.480 1092.500 870.280 ;
        RECT 149.620 853.280 594.720 858.480 ;
        RECT 149.620 810.480 1092.500 853.280 ;
        RECT 149.620 805.280 594.720 810.480 ;
        RECT 149.620 793.480 1092.500 805.280 ;
        RECT 237.800 788.280 421.560 793.480 ;
        RECT 149.620 745.480 1092.500 788.280 ;
        RECT 237.800 740.280 421.560 745.480 ;
        RECT 149.620 728.480 1092.500 740.280 ;
        RECT 237.800 723.280 421.560 728.480 ;
        RECT 149.620 680.480 1092.500 723.280 ;
        RECT 237.800 675.280 421.560 680.480 ;
        RECT 149.620 663.480 1092.500 675.280 ;
        RECT 149.620 658.280 594.720 663.480 ;
        RECT 149.620 615.480 1092.500 658.280 ;
        RECT 237.800 610.280 574.600 615.480 ;
        RECT 149.620 598.480 1092.500 610.280 ;
        RECT 149.620 593.280 594.720 598.480 ;
        RECT 149.620 550.480 1092.500 593.280 ;
        RECT 149.620 545.280 594.720 550.480 ;
        RECT 149.620 533.480 1092.500 545.280 ;
        RECT 149.620 527.900 1092.500 528.280 ;
        RECT 614.720 522.700 1092.500 527.900 ;
        RECT 149.620 485.480 1092.500 522.700 ;
        RECT 149.620 468.480 1092.500 480.280 ;
        RECT 149.620 463.280 594.720 468.480 ;
        RECT 149.620 420.480 1092.500 463.280 ;
        RECT 149.620 415.280 594.720 420.480 ;
        RECT 149.620 403.480 1092.500 415.280 ;
        RECT 149.620 398.280 594.720 403.480 ;
        RECT 149.620 355.480 1092.500 398.280 ;
        RECT 149.620 350.280 594.720 355.480 ;
        RECT 149.620 338.480 1092.500 350.280 ;
        RECT 149.620 333.280 594.720 338.480 ;
        RECT 149.620 290.480 1092.500 333.280 ;
        RECT 149.620 285.280 594.720 290.480 ;
        RECT 149.620 273.480 1092.500 285.280 ;
        RECT 237.800 268.280 421.560 273.480 ;
        RECT 149.620 225.480 1092.500 268.280 ;
        RECT 149.620 220.280 594.720 225.480 ;
        RECT 149.620 208.480 1092.500 220.280 ;
        RECT 237.800 203.280 464.930 208.480 ;
        RECT 149.620 160.480 1092.500 203.280 ;
        RECT 237.800 155.280 574.600 160.480 ;
        RECT 149.620 143.480 1092.500 155.280 ;
        RECT 149.620 138.280 594.720 143.480 ;
        RECT 149.620 99.980 1092.500 138.280 ;
  END
END signal_generator
END LIBRARY

