VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO designs_wrapper
  CLASS BLOCK ;
  FOREIGN designs_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2000.000 BY 900.000 ;
  PIN i_clock
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 448.840 4.000 449.440 ;
    END
  END i_clock
  PIN i_enable
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 788.840 4.000 789.440 ;
    END
  END i_enable
  PIN i_freq_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 516.840 4.000 517.440 ;
    END
  END i_freq_sel[0]
  PIN i_freq_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 584.840 4.000 585.440 ;
    END
  END i_freq_sel[1]
  PIN i_freq_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 652.840 4.000 653.440 ;
    END
  END i_freq_sel[2]
  PIN i_freq_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 720.840 4.000 721.440 ;
    END
  END i_freq_sel[3]
  PIN i_signal_sel
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 856.840 4.000 857.440 ;
    END
  END i_signal_sel
  PIN i_test
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.840 4.000 381.440 ;
    END
  END i_test
  PIN i_wb_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 719.530 0.000 719.810 4.000 ;
    END
  END i_wb_addr[0]
  PIN i_wb_addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 526.330 0.000 526.610 4.000 ;
    END
  END i_wb_addr[10]
  PIN i_wb_addr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 507.010 0.000 507.290 4.000 ;
    END
  END i_wb_addr[11]
  PIN i_wb_addr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 487.690 0.000 487.970 4.000 ;
    END
  END i_wb_addr[12]
  PIN i_wb_addr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 468.370 0.000 468.650 4.000 ;
    END
  END i_wb_addr[13]
  PIN i_wb_addr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 449.050 0.000 449.330 4.000 ;
    END
  END i_wb_addr[14]
  PIN i_wb_addr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 429.730 0.000 430.010 4.000 ;
    END
  END i_wb_addr[15]
  PIN i_wb_addr[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 410.410 0.000 410.690 4.000 ;
    END
  END i_wb_addr[16]
  PIN i_wb_addr[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 391.090 0.000 391.370 4.000 ;
    END
  END i_wb_addr[17]
  PIN i_wb_addr[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 371.770 0.000 372.050 4.000 ;
    END
  END i_wb_addr[18]
  PIN i_wb_addr[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 352.450 0.000 352.730 4.000 ;
    END
  END i_wb_addr[19]
  PIN i_wb_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 700.210 0.000 700.490 4.000 ;
    END
  END i_wb_addr[1]
  PIN i_wb_addr[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 333.130 0.000 333.410 4.000 ;
    END
  END i_wb_addr[20]
  PIN i_wb_addr[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 313.810 0.000 314.090 4.000 ;
    END
  END i_wb_addr[21]
  PIN i_wb_addr[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 294.490 0.000 294.770 4.000 ;
    END
  END i_wb_addr[22]
  PIN i_wb_addr[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 275.170 0.000 275.450 4.000 ;
    END
  END i_wb_addr[23]
  PIN i_wb_addr[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 255.850 0.000 256.130 4.000 ;
    END
  END i_wb_addr[24]
  PIN i_wb_addr[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 236.530 0.000 236.810 4.000 ;
    END
  END i_wb_addr[25]
  PIN i_wb_addr[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 217.210 0.000 217.490 4.000 ;
    END
  END i_wb_addr[26]
  PIN i_wb_addr[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 197.890 0.000 198.170 4.000 ;
    END
  END i_wb_addr[27]
  PIN i_wb_addr[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 178.570 0.000 178.850 4.000 ;
    END
  END i_wb_addr[28]
  PIN i_wb_addr[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 159.250 0.000 159.530 4.000 ;
    END
  END i_wb_addr[29]
  PIN i_wb_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 680.890 0.000 681.170 4.000 ;
    END
  END i_wb_addr[2]
  PIN i_wb_addr[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 139.930 0.000 140.210 4.000 ;
    END
  END i_wb_addr[30]
  PIN i_wb_addr[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 120.610 0.000 120.890 4.000 ;
    END
  END i_wb_addr[31]
  PIN i_wb_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 661.570 0.000 661.850 4.000 ;
    END
  END i_wb_addr[3]
  PIN i_wb_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 642.250 0.000 642.530 4.000 ;
    END
  END i_wb_addr[4]
  PIN i_wb_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 622.930 0.000 623.210 4.000 ;
    END
  END i_wb_addr[5]
  PIN i_wb_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 603.610 0.000 603.890 4.000 ;
    END
  END i_wb_addr[6]
  PIN i_wb_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 584.290 0.000 584.570 4.000 ;
    END
  END i_wb_addr[7]
  PIN i_wb_addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 564.970 0.000 565.250 4.000 ;
    END
  END i_wb_addr[8]
  PIN i_wb_addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 545.650 0.000 545.930 4.000 ;
    END
  END i_wb_addr[9]
  PIN i_wb_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 24.010 0.000 24.290 4.000 ;
    END
  END i_wb_clk
  PIN i_wb_cyc
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 62.650 0.000 62.930 4.000 ;
    END
  END i_wb_cyc
  PIN i_wb_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 1337.770 0.000 1338.050 4.000 ;
    END
  END i_wb_data[0]
  PIN i_wb_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1144.570 0.000 1144.850 4.000 ;
    END
  END i_wb_data[10]
  PIN i_wb_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1125.250 0.000 1125.530 4.000 ;
    END
  END i_wb_data[11]
  PIN i_wb_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1105.930 0.000 1106.210 4.000 ;
    END
  END i_wb_data[12]
  PIN i_wb_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1086.610 0.000 1086.890 4.000 ;
    END
  END i_wb_data[13]
  PIN i_wb_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1067.290 0.000 1067.570 4.000 ;
    END
  END i_wb_data[14]
  PIN i_wb_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1047.970 0.000 1048.250 4.000 ;
    END
  END i_wb_data[15]
  PIN i_wb_data[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1028.650 0.000 1028.930 4.000 ;
    END
  END i_wb_data[16]
  PIN i_wb_data[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1009.330 0.000 1009.610 4.000 ;
    END
  END i_wb_data[17]
  PIN i_wb_data[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 990.010 0.000 990.290 4.000 ;
    END
  END i_wb_data[18]
  PIN i_wb_data[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 970.690 0.000 970.970 4.000 ;
    END
  END i_wb_data[19]
  PIN i_wb_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 1318.450 0.000 1318.730 4.000 ;
    END
  END i_wb_data[1]
  PIN i_wb_data[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 951.370 0.000 951.650 4.000 ;
    END
  END i_wb_data[20]
  PIN i_wb_data[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 932.050 0.000 932.330 4.000 ;
    END
  END i_wb_data[21]
  PIN i_wb_data[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 912.730 0.000 913.010 4.000 ;
    END
  END i_wb_data[22]
  PIN i_wb_data[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 893.410 0.000 893.690 4.000 ;
    END
  END i_wb_data[23]
  PIN i_wb_data[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 874.090 0.000 874.370 4.000 ;
    END
  END i_wb_data[24]
  PIN i_wb_data[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 854.770 0.000 855.050 4.000 ;
    END
  END i_wb_data[25]
  PIN i_wb_data[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 835.450 0.000 835.730 4.000 ;
    END
  END i_wb_data[26]
  PIN i_wb_data[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 816.130 0.000 816.410 4.000 ;
    END
  END i_wb_data[27]
  PIN i_wb_data[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 796.810 0.000 797.090 4.000 ;
    END
  END i_wb_data[28]
  PIN i_wb_data[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 777.490 0.000 777.770 4.000 ;
    END
  END i_wb_data[29]
  PIN i_wb_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 1299.130 0.000 1299.410 4.000 ;
    END
  END i_wb_data[2]
  PIN i_wb_data[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 758.170 0.000 758.450 4.000 ;
    END
  END i_wb_data[30]
  PIN i_wb_data[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 738.850 0.000 739.130 4.000 ;
    END
  END i_wb_data[31]
  PIN i_wb_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 1279.810 0.000 1280.090 4.000 ;
    END
  END i_wb_data[3]
  PIN i_wb_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1260.490 0.000 1260.770 4.000 ;
    END
  END i_wb_data[4]
  PIN i_wb_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1241.170 0.000 1241.450 4.000 ;
    END
  END i_wb_data[5]
  PIN i_wb_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1221.850 0.000 1222.130 4.000 ;
    END
  END i_wb_data[6]
  PIN i_wb_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1202.530 0.000 1202.810 4.000 ;
    END
  END i_wb_data[7]
  PIN i_wb_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1183.210 0.000 1183.490 4.000 ;
    END
  END i_wb_data[8]
  PIN i_wb_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1163.890 0.000 1164.170 4.000 ;
    END
  END i_wb_data[9]
  PIN i_wb_rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 43.330 0.000 43.610 4.000 ;
    END
  END i_wb_rst
  PIN i_wb_stb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 81.970 0.000 82.250 4.000 ;
    END
  END i_wb_stb
  PIN i_wb_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 101.290 0.000 101.570 4.000 ;
    END
  END i_wb_we
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 873.160 2000.000 873.760 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 546.760 2000.000 547.360 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 514.120 2000.000 514.720 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 481.480 2000.000 482.080 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 448.840 2000.000 449.440 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 416.200 2000.000 416.800 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 383.560 2000.000 384.160 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 350.920 2000.000 351.520 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 318.280 2000.000 318.880 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 285.640 2000.000 286.240 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 253.000 2000.000 253.600 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 840.520 2000.000 841.120 ;
    END
  END io_oeb[1]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 807.880 2000.000 808.480 ;
    END
  END io_oeb[2]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 775.240 2000.000 775.840 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 742.600 2000.000 743.200 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 709.960 2000.000 710.560 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 677.320 2000.000 677.920 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 644.680 2000.000 645.280 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 612.040 2000.000 612.640 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 579.400 2000.000 580.000 ;
    END
  END io_oeb[9]
  PIN o_ADC_frame
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 1996.000 57.160 2000.000 57.760 ;
    END
  END o_ADC_frame
  PIN o_control_signal
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 1996.000 220.360 2000.000 220.960 ;
    END
  END o_control_signal
  PIN o_phi_l1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 1996.000 89.800 2000.000 90.400 ;
    END
  END o_phi_l1
  PIN o_phi_l2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 1996.000 122.440 2000.000 123.040 ;
    END
  END o_phi_l2
  PIN o_phi_p
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 1996.000 155.080 2000.000 155.680 ;
    END
  END o_phi_p
  PIN o_phi_r
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 1996.000 187.720 2000.000 188.320 ;
    END
  END o_phi_r
  PIN o_pixel_flag
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 1996.000 24.520 2000.000 25.120 ;
    END
  END o_pixel_flag
  PIN o_test[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END o_test[0]
  PIN o_test[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END o_test[1]
  PIN o_test[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END o_test[2]
  PIN o_test[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.840 4.000 245.440 ;
    END
  END o_test[3]
  PIN o_test[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.840 4.000 313.440 ;
    END
  END o_test[4]
  PIN o_wb_ack
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1357.090 0.000 1357.370 4.000 ;
    END
  END o_wb_ack
  PIN o_wb_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1975.330 0.000 1975.610 4.000 ;
    END
  END o_wb_data[0]
  PIN o_wb_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1782.130 0.000 1782.410 4.000 ;
    END
  END o_wb_data[10]
  PIN o_wb_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1762.810 0.000 1763.090 4.000 ;
    END
  END o_wb_data[11]
  PIN o_wb_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1743.490 0.000 1743.770 4.000 ;
    END
  END o_wb_data[12]
  PIN o_wb_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1724.170 0.000 1724.450 4.000 ;
    END
  END o_wb_data[13]
  PIN o_wb_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1704.850 0.000 1705.130 4.000 ;
    END
  END o_wb_data[14]
  PIN o_wb_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1685.530 0.000 1685.810 4.000 ;
    END
  END o_wb_data[15]
  PIN o_wb_data[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1666.210 0.000 1666.490 4.000 ;
    END
  END o_wb_data[16]
  PIN o_wb_data[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1646.890 0.000 1647.170 4.000 ;
    END
  END o_wb_data[17]
  PIN o_wb_data[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1627.570 0.000 1627.850 4.000 ;
    END
  END o_wb_data[18]
  PIN o_wb_data[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1608.250 0.000 1608.530 4.000 ;
    END
  END o_wb_data[19]
  PIN o_wb_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1956.010 0.000 1956.290 4.000 ;
    END
  END o_wb_data[1]
  PIN o_wb_data[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1588.930 0.000 1589.210 4.000 ;
    END
  END o_wb_data[20]
  PIN o_wb_data[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1569.610 0.000 1569.890 4.000 ;
    END
  END o_wb_data[21]
  PIN o_wb_data[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1550.290 0.000 1550.570 4.000 ;
    END
  END o_wb_data[22]
  PIN o_wb_data[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1530.970 0.000 1531.250 4.000 ;
    END
  END o_wb_data[23]
  PIN o_wb_data[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1511.650 0.000 1511.930 4.000 ;
    END
  END o_wb_data[24]
  PIN o_wb_data[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1492.330 0.000 1492.610 4.000 ;
    END
  END o_wb_data[25]
  PIN o_wb_data[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1473.010 0.000 1473.290 4.000 ;
    END
  END o_wb_data[26]
  PIN o_wb_data[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1453.690 0.000 1453.970 4.000 ;
    END
  END o_wb_data[27]
  PIN o_wb_data[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1434.370 0.000 1434.650 4.000 ;
    END
  END o_wb_data[28]
  PIN o_wb_data[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1415.050 0.000 1415.330 4.000 ;
    END
  END o_wb_data[29]
  PIN o_wb_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1936.690 0.000 1936.970 4.000 ;
    END
  END o_wb_data[2]
  PIN o_wb_data[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1395.730 0.000 1396.010 4.000 ;
    END
  END o_wb_data[30]
  PIN o_wb_data[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1376.410 0.000 1376.690 4.000 ;
    END
  END o_wb_data[31]
  PIN o_wb_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1917.370 0.000 1917.650 4.000 ;
    END
  END o_wb_data[3]
  PIN o_wb_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1898.050 0.000 1898.330 4.000 ;
    END
  END o_wb_data[4]
  PIN o_wb_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1878.730 0.000 1879.010 4.000 ;
    END
  END o_wb_data[5]
  PIN o_wb_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1859.410 0.000 1859.690 4.000 ;
    END
  END o_wb_data[6]
  PIN o_wb_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1840.090 0.000 1840.370 4.000 ;
    END
  END o_wb_data[7]
  PIN o_wb_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1820.770 0.000 1821.050 4.000 ;
    END
  END o_wb_data[8]
  PIN o_wb_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1801.450 0.000 1801.730 4.000 ;
    END
  END o_wb_data[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1557.040 10.640 1558.640 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1710.640 10.640 1712.240 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1864.240 10.640 1865.840 886.960 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1633.840 10.640 1635.440 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1787.440 10.640 1789.040 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1941.040 10.640 1942.640 886.960 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1994.100 886.805 ;
      LAYER met1 ;
        RECT 4.670 8.880 1994.100 886.960 ;
      LAYER met2 ;
        RECT 4.690 4.280 1992.630 886.905 ;
        RECT 4.690 3.670 23.730 4.280 ;
        RECT 24.570 3.670 43.050 4.280 ;
        RECT 43.890 3.670 62.370 4.280 ;
        RECT 63.210 3.670 81.690 4.280 ;
        RECT 82.530 3.670 101.010 4.280 ;
        RECT 101.850 3.670 120.330 4.280 ;
        RECT 121.170 3.670 139.650 4.280 ;
        RECT 140.490 3.670 158.970 4.280 ;
        RECT 159.810 3.670 178.290 4.280 ;
        RECT 179.130 3.670 197.610 4.280 ;
        RECT 198.450 3.670 216.930 4.280 ;
        RECT 217.770 3.670 236.250 4.280 ;
        RECT 237.090 3.670 255.570 4.280 ;
        RECT 256.410 3.670 274.890 4.280 ;
        RECT 275.730 3.670 294.210 4.280 ;
        RECT 295.050 3.670 313.530 4.280 ;
        RECT 314.370 3.670 332.850 4.280 ;
        RECT 333.690 3.670 352.170 4.280 ;
        RECT 353.010 3.670 371.490 4.280 ;
        RECT 372.330 3.670 390.810 4.280 ;
        RECT 391.650 3.670 410.130 4.280 ;
        RECT 410.970 3.670 429.450 4.280 ;
        RECT 430.290 3.670 448.770 4.280 ;
        RECT 449.610 3.670 468.090 4.280 ;
        RECT 468.930 3.670 487.410 4.280 ;
        RECT 488.250 3.670 506.730 4.280 ;
        RECT 507.570 3.670 526.050 4.280 ;
        RECT 526.890 3.670 545.370 4.280 ;
        RECT 546.210 3.670 564.690 4.280 ;
        RECT 565.530 3.670 584.010 4.280 ;
        RECT 584.850 3.670 603.330 4.280 ;
        RECT 604.170 3.670 622.650 4.280 ;
        RECT 623.490 3.670 641.970 4.280 ;
        RECT 642.810 3.670 661.290 4.280 ;
        RECT 662.130 3.670 680.610 4.280 ;
        RECT 681.450 3.670 699.930 4.280 ;
        RECT 700.770 3.670 719.250 4.280 ;
        RECT 720.090 3.670 738.570 4.280 ;
        RECT 739.410 3.670 757.890 4.280 ;
        RECT 758.730 3.670 777.210 4.280 ;
        RECT 778.050 3.670 796.530 4.280 ;
        RECT 797.370 3.670 815.850 4.280 ;
        RECT 816.690 3.670 835.170 4.280 ;
        RECT 836.010 3.670 854.490 4.280 ;
        RECT 855.330 3.670 873.810 4.280 ;
        RECT 874.650 3.670 893.130 4.280 ;
        RECT 893.970 3.670 912.450 4.280 ;
        RECT 913.290 3.670 931.770 4.280 ;
        RECT 932.610 3.670 951.090 4.280 ;
        RECT 951.930 3.670 970.410 4.280 ;
        RECT 971.250 3.670 989.730 4.280 ;
        RECT 990.570 3.670 1009.050 4.280 ;
        RECT 1009.890 3.670 1028.370 4.280 ;
        RECT 1029.210 3.670 1047.690 4.280 ;
        RECT 1048.530 3.670 1067.010 4.280 ;
        RECT 1067.850 3.670 1086.330 4.280 ;
        RECT 1087.170 3.670 1105.650 4.280 ;
        RECT 1106.490 3.670 1124.970 4.280 ;
        RECT 1125.810 3.670 1144.290 4.280 ;
        RECT 1145.130 3.670 1163.610 4.280 ;
        RECT 1164.450 3.670 1182.930 4.280 ;
        RECT 1183.770 3.670 1202.250 4.280 ;
        RECT 1203.090 3.670 1221.570 4.280 ;
        RECT 1222.410 3.670 1240.890 4.280 ;
        RECT 1241.730 3.670 1260.210 4.280 ;
        RECT 1261.050 3.670 1279.530 4.280 ;
        RECT 1280.370 3.670 1298.850 4.280 ;
        RECT 1299.690 3.670 1318.170 4.280 ;
        RECT 1319.010 3.670 1337.490 4.280 ;
        RECT 1338.330 3.670 1356.810 4.280 ;
        RECT 1357.650 3.670 1376.130 4.280 ;
        RECT 1376.970 3.670 1395.450 4.280 ;
        RECT 1396.290 3.670 1414.770 4.280 ;
        RECT 1415.610 3.670 1434.090 4.280 ;
        RECT 1434.930 3.670 1453.410 4.280 ;
        RECT 1454.250 3.670 1472.730 4.280 ;
        RECT 1473.570 3.670 1492.050 4.280 ;
        RECT 1492.890 3.670 1511.370 4.280 ;
        RECT 1512.210 3.670 1530.690 4.280 ;
        RECT 1531.530 3.670 1550.010 4.280 ;
        RECT 1550.850 3.670 1569.330 4.280 ;
        RECT 1570.170 3.670 1588.650 4.280 ;
        RECT 1589.490 3.670 1607.970 4.280 ;
        RECT 1608.810 3.670 1627.290 4.280 ;
        RECT 1628.130 3.670 1646.610 4.280 ;
        RECT 1647.450 3.670 1665.930 4.280 ;
        RECT 1666.770 3.670 1685.250 4.280 ;
        RECT 1686.090 3.670 1704.570 4.280 ;
        RECT 1705.410 3.670 1723.890 4.280 ;
        RECT 1724.730 3.670 1743.210 4.280 ;
        RECT 1744.050 3.670 1762.530 4.280 ;
        RECT 1763.370 3.670 1781.850 4.280 ;
        RECT 1782.690 3.670 1801.170 4.280 ;
        RECT 1802.010 3.670 1820.490 4.280 ;
        RECT 1821.330 3.670 1839.810 4.280 ;
        RECT 1840.650 3.670 1859.130 4.280 ;
        RECT 1859.970 3.670 1878.450 4.280 ;
        RECT 1879.290 3.670 1897.770 4.280 ;
        RECT 1898.610 3.670 1917.090 4.280 ;
        RECT 1917.930 3.670 1936.410 4.280 ;
        RECT 1937.250 3.670 1955.730 4.280 ;
        RECT 1956.570 3.670 1975.050 4.280 ;
        RECT 1975.890 3.670 1992.630 4.280 ;
      LAYER met3 ;
        RECT 4.000 874.160 1996.000 886.885 ;
        RECT 4.000 872.760 1995.600 874.160 ;
        RECT 4.000 857.840 1996.000 872.760 ;
        RECT 4.400 856.440 1996.000 857.840 ;
        RECT 4.000 841.520 1996.000 856.440 ;
        RECT 4.000 840.120 1995.600 841.520 ;
        RECT 4.000 808.880 1996.000 840.120 ;
        RECT 4.000 807.480 1995.600 808.880 ;
        RECT 4.000 789.840 1996.000 807.480 ;
        RECT 4.400 788.440 1996.000 789.840 ;
        RECT 4.000 776.240 1996.000 788.440 ;
        RECT 4.000 774.840 1995.600 776.240 ;
        RECT 4.000 743.600 1996.000 774.840 ;
        RECT 4.000 742.200 1995.600 743.600 ;
        RECT 4.000 721.840 1996.000 742.200 ;
        RECT 4.400 720.440 1996.000 721.840 ;
        RECT 4.000 710.960 1996.000 720.440 ;
        RECT 4.000 709.560 1995.600 710.960 ;
        RECT 4.000 678.320 1996.000 709.560 ;
        RECT 4.000 676.920 1995.600 678.320 ;
        RECT 4.000 653.840 1996.000 676.920 ;
        RECT 4.400 652.440 1996.000 653.840 ;
        RECT 4.000 645.680 1996.000 652.440 ;
        RECT 4.000 644.280 1995.600 645.680 ;
        RECT 4.000 613.040 1996.000 644.280 ;
        RECT 4.000 611.640 1995.600 613.040 ;
        RECT 4.000 585.840 1996.000 611.640 ;
        RECT 4.400 584.440 1996.000 585.840 ;
        RECT 4.000 580.400 1996.000 584.440 ;
        RECT 4.000 579.000 1995.600 580.400 ;
        RECT 4.000 547.760 1996.000 579.000 ;
        RECT 4.000 546.360 1995.600 547.760 ;
        RECT 4.000 517.840 1996.000 546.360 ;
        RECT 4.400 516.440 1996.000 517.840 ;
        RECT 4.000 515.120 1996.000 516.440 ;
        RECT 4.000 513.720 1995.600 515.120 ;
        RECT 4.000 482.480 1996.000 513.720 ;
        RECT 4.000 481.080 1995.600 482.480 ;
        RECT 4.000 449.840 1996.000 481.080 ;
        RECT 4.400 448.440 1995.600 449.840 ;
        RECT 4.000 417.200 1996.000 448.440 ;
        RECT 4.000 415.800 1995.600 417.200 ;
        RECT 4.000 384.560 1996.000 415.800 ;
        RECT 4.000 383.160 1995.600 384.560 ;
        RECT 4.000 381.840 1996.000 383.160 ;
        RECT 4.400 380.440 1996.000 381.840 ;
        RECT 4.000 351.920 1996.000 380.440 ;
        RECT 4.000 350.520 1995.600 351.920 ;
        RECT 4.000 319.280 1996.000 350.520 ;
        RECT 4.000 317.880 1995.600 319.280 ;
        RECT 4.000 313.840 1996.000 317.880 ;
        RECT 4.400 312.440 1996.000 313.840 ;
        RECT 4.000 286.640 1996.000 312.440 ;
        RECT 4.000 285.240 1995.600 286.640 ;
        RECT 4.000 254.000 1996.000 285.240 ;
        RECT 4.000 252.600 1995.600 254.000 ;
        RECT 4.000 245.840 1996.000 252.600 ;
        RECT 4.400 244.440 1996.000 245.840 ;
        RECT 4.000 221.360 1996.000 244.440 ;
        RECT 4.000 219.960 1995.600 221.360 ;
        RECT 4.000 188.720 1996.000 219.960 ;
        RECT 4.000 187.320 1995.600 188.720 ;
        RECT 4.000 177.840 1996.000 187.320 ;
        RECT 4.400 176.440 1996.000 177.840 ;
        RECT 4.000 156.080 1996.000 176.440 ;
        RECT 4.000 154.680 1995.600 156.080 ;
        RECT 4.000 123.440 1996.000 154.680 ;
        RECT 4.000 122.040 1995.600 123.440 ;
        RECT 4.000 109.840 1996.000 122.040 ;
        RECT 4.400 108.440 1996.000 109.840 ;
        RECT 4.000 90.800 1996.000 108.440 ;
        RECT 4.000 89.400 1995.600 90.800 ;
        RECT 4.000 58.160 1996.000 89.400 ;
        RECT 4.000 56.760 1995.600 58.160 ;
        RECT 4.000 41.840 1996.000 56.760 ;
        RECT 4.400 40.440 1996.000 41.840 ;
        RECT 4.000 25.520 1996.000 40.440 ;
        RECT 4.000 24.120 1995.600 25.520 ;
        RECT 4.000 10.715 1996.000 24.120 ;
  END
END designs_wrapper
END LIBRARY

